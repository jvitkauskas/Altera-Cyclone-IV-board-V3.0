module half_adder(
    A,					//����ѡ���ַ�ɿ��ؾ�����0�����£�1��δ����
	B,					//����ѡ���ַ�ɿ��ؾ�����0�����£�1��δ����
	
	S,					//�����0��������1��Ϩ��
	C					//�����0��������1��Ϩ��
    );
input			A;			//����˿�
input			B;			//����˿�

output		S;			//����˿�
output		C;			//����˿�

assign S = A ^ B;				//ֱ�Ӹ�ֵ�����
assign C = A & B;			//ֱ�Ӹ�ֵ����

endmodule
