��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�+����Rq�����������+�nS�U�F7&���S����"�M ��U���@�˴�5��.� -;P�~�oa|
)k���BЖ�@�o�v�4ߘ<��4�l��D�4Ak���-.b���mC*��D�i�M%��%�k�~&ʳ��0!����nY�qe��3��ck����o��z"��,f�ը��%$���|�;+#�0f�UhOǃ��2刑�Lc�����|��|����Q��Ol�pf��\�4Y�
A�Y�a@��qnNAz�pד��ݮiF�?��'~&{�X�v����H�	���Gʲ���dӤ�>v�� ���K�B�x��X�[#s��W�V��.��f$�n���:Qn��24"M��<48�}[�� �(�5��t�L�6����ئe3Xa�|=�X$nD�H"ď�Vl��⼞=��5��n�Q���6;#٬"I�L���P����/P=�}�㟂���C���?�ZI�r�	5��]%���ē�2FTC�Sh��Ds]鉬�@�0:�?"ܮAۙ�>���?��i+c��$�vf�:��P����LX�Z��+�'��Y�}�G��)��q��ʋ�X�]���ۅЅ�aڴG��i����(ް?	�P9���y�
�����E==6�iS��=م�gU����!��8�د�§���g��d���B�Rx%��E}��8�!-�U��@=�R ��s�/�ǥ�;,'�f��|�<�\W�21u�a���{-��������k�����@b��G�9SK{[O��Y��7�vb���yS�����	�63ǲ�Sr�,B�/�t�(��� bc";W���"-�����?�1\�ؤ'

`�x��4Q.�H����E�l���5��S���kd1��{+Hڔ�խ8�|$�������؄+����)���gn��+砯y���>3T��Xw5ӗ<,�C���   ̰�78ys
7�s�m�MO���_���t�3���d���*�۱�)!܃�9��-�J���.��qkT�*)�
0�Fx����t�g#@p��s���(��ܐ�q��U)ײ�Zƚś�!����qp� }�̚ޒ��	�v4V���t"��V�fn��΂��^� !��!G����Db�sU���9����n�)��n�oŠvs�m]��ʐ��ǌ���8$��
M5�I8G��	����EG��.N6���i��5pX�\��Z���>s�EY��Wo��OQ7�π����`�|�B6_V��39���b�b��U��Zn�8��4�&�^�3��.�ߊ&��B�g`��L�+4��m�	Ɛ�=���u�JR�)��
�%	���Y����v���h<�ŝA��OU�9��x'���N��^[#�k4+��4�]M\�$
��!�&�{�Y.KY���̈́��'5B$(��;�6�.:+U��;Y�3�6ݱT����T����~F4������-`����M��s�t ���Z���-����,+�ج�pYkk�x��&��Y,����ZA��vז�&��ý����Oʺ���"}@B\�x�sV<��j�VӴ�'�礣\գ>58^��z�����9���k�G��ɣ�У^�x_��]\Z����ֈ�S��5Pf)����H���U
$��-��t�!���^4?�����~e2��@�a��
Ȑ�+��)��_�T·R����ln���,PꪶX��?{fo�b^;퇈E�??�c� �u���d�\i.R����6d�8�IZȗ�@ȹIc�"�9�nG�崕^P���,GF�Ð�s"�\�7�@��ޯ�F�$���eb=`�Al�^{�l�#SL�7��G§����ri�ha�J�Ē��6�*m=�WNKÐZ�(��u��V8<a�M���|I��r�Q�ah�[�{^e��ָ�w\~bI��ĴWӺΡ��D�0���_��_������ǷS�)�K���A���(��i��"��'�A��3s��D�64�hڷ׸���h�A�,;t/AhP�A�:T�"{�����?�"c���8��e�,޸��]�:6�*e0�>�j]�cǩ�2Ns��n'c>��q �T &7�d��s���z�$�a��{ކE�.���ORj�փ�}_C]�e�gO7}����D���H��|�*'!�$J٬/��Բ@p��x5}���7�������q:rIWo���loKTЁ@采oB�l��lp����B|ת��ӀP_޾p��U}��Bmp�v&�ʟ���$�1�����Ɗ������BQ�U�*��������	5�U�׵a�"(JH��@�rsoh	oA�x`���.��K��k3��1m7A���|�U��)��z�]�ԉR�+�[<lP�aze!׳��}|�P���:S�jɟ5�cO�Q��]�u}�k�T&iw��~`�z!r��~A�C�����9}?��t�s��>$I���$Ի֖c�ӟ�Nv�x���#�Չ���{=�2��9z�C�J�9�s���Ϭ�%6�_�2�{��<�?�a&dҘ|����"�x]8Z�>:��"�F��2 э-a���9)�գD������������%X��ϩ�����CI���%�k�!��g@ ���ǽN� &�kV��O:��C4P�j��=]�V�\zX���O	��b��CҴ�H�8��|�]N]���vJ�ɲ[ H��H"D�J��h��t�gJ��$�nmE�>���Q�l���^��` ɮ�l�4o�(v���s�q�76��q#�6�4�Kw�'7�ZHoht�`?UN���M�	M<�7ƃ�n�=�6=u���=���j����(z<>���/y�?v����О�$��m�'�G�M�]:-D��}��uza$����_b3ӗςE����T�
G�֜�Rb�5���^w���_j��k
�i�V��.l#2�e�&N�����b)����g�ܘ���L(�$��(M$>��q��3���x8�DC��S�u�4�Q�Ġ�SFȵFp��l.%�ȯz���y����:�|1�vUB9�jo;T-�<�s3�\br@;q6/�#{����T��xV�L#�#��_��
ܺ�f�@���{�(���P��cU�]�ǭ2�[� ���g��MN�n��c��ꔃW�[`�I@j��^�PՁU��.�$��:�m+�� ��� ՘��S�0��E�UDLd�	eqQ;VL+X�7���{d��Qo�׏��h�`/
�cc�9ŋKs�r�߻��x��%*�>޹J��C��\�`C1OI���;ݛ ������i
��45P���>ť�8�S�@ 0�Ƅ.�1E�uȁ}���Y���Gc��/[w�6*[��D�o���o��f>�w�"����J>�����@@ADN|�3��d��'0<����kE?#��dV; �o�Q�N�Xn1��S�)���ZuT�� "ka�_���2;1�
��No��?D ���t�B�V��ƪ��wln�:V�(���dHW%u��<@�S��A��l�8];Qa�L�9$^%� �i0,���u\E�'�*�ț�u���%=�
u�O�p�C�=��uؿ�z�x+���������`����)c�X��l��S��v�k�Λ�\"�r��@��k�]��/@��3a��' Bݘ|�DZ���a�ֹ�Z����h����X	���kV�5$ڋ\z��͉��;����0E�ƛ��j'Y�������7$�Y�Sܓ�X��vV2�F�2ί�XﱂB��
=�N��>Ӓ�)��N���f��X:�WQ^3��t����jO��������ѽ�������^oSc�m�g�ی;ű�!qG��agy�D�Y!s1��_Jů?k�y�����e=��	|)�N��\Y���R�~Y}�I�WwUh�������� ���
�jv,j`����f�Y�c�⛺%�JW��pLn?�ʢ����C��F�����;Zf��#��ʔ46Ǐ {�څ�Q��m�����pP�g�W��-�Bx�c���&ʈ�鷥�e���OG��@�sv�n =�z�bBj��1C��.̩�)��@d���,�O��͍h0�=�^��R����nq ]�m�6e�f�H�`�߂�����+�i��7���k��S��=~ϝ	���"$����b/�����r+X#�Lm�l&�,�����.kDL+;�n��; �$�h	cA(�@x6�X;�͞s\�E�$Aj�Vk�a
M�O���?�[R�	!�Kpp����k���40@e"u��E����L�G�5;��Z��s�����w��q�ȭ�翣���h*�ے:���
�c�#+�⣩�
�7��1]���l�,� z(�<�[��V�)5FĿH;�vD:㝖�F�)s@@�U4q{ |�?1k�s�=�\^E���Bӓ/��]�nr�#�.�����r��� �jD	-^� �������rNG�"y�{����^���B��*|z����b�]/S�.Y%����ܢ\�ú���K���5����߅(D�u� ¹f#'Y6����I��#�)x�c�*)o��E0\*�R5*���U����Q3#
Ҹ��\۶��9���"=�Li��ki�0�m���c���p̊�("kG"t3�oNZ,�)��݆.��C�אv��/�W�W����U��\��	�G�"sѡ��(���� ���������^1$?�Ί�X��t�s�h�!�;��p\�hU|��7�Я������t����I��s)�@�*�M���r9�y�t:�c���ߦ��6 �L�}�Z�n��[��-*�M����ߐ��
yPq�H!��H������RX*g�������`{���&�&6�ULt�)��g@�^g�6�Ī2g��BcC����|�j��bvz�6��t@J���>��T��Hy#�|�͐��#�`�˂8Y��������i���-�ï��^<���z�Y�AL���d�F�x�Z�D9�+cdE��M ���gcu��Gu.�>��$Q|���f�Άٖ@[S�6ޟp0d�LZ�n�|G������4=�h��*�{��8���-�_v��C���Ş}4H�V�Vp&d�M.k:hFY�2 �ܽM��W�':Y����Ӵf�oĐ��S���ۻ�NM�!�T\D�.Rk�
Wu�TZ�"T��JMKSՀ��iv�pB��n�-<��.0H�u)M��_�J3zg ��n�R��Cuu�qf.�ƿ���|��t;w�ﭨ��_���d����}[����ư7�8sf�w$�������O_����1��H��%+��>a���#��ӽ��m�F��l>�[ɾ������Z������0�	���]���(Y@�w�݆Ǩ<��q�(�5�s�ej�I���&�v]�+b���*��>��X�2*c���E����D����7�r ���MA�j ��p����3��_xAl���4/��2�(�
?JB �H(���|񧿙��O��3��-���m�<v��sD���@�f��&�(
�I<#7����ޔ��u���:�G�����j;��E�����[�� ��I�������1JDI�nq�LQ,���b0��,J@5�E � ��`@C<��,Z�f������C�7��1�k��^x�z�慍���5����)\y���� ���-Z�z4i��\j�SN�d#͜�.ܛ��Yq��|x����>�����,wN>���0����9 �x���C�Wd�� q���$)zpxV͡-�X*�Zif!���EUţ9�g�?��9���H*G��C}����b�����������i��s)������V�⡦�m@��l�,0{��]�]��;<ՌtYq-p`��F��#�K�m�D�����w��
4�4�<�7f\78��S�BZ�crw@M@��co�ۿ��Qqe�����QO<��J�Q�?�[���_�&�r �]߹b�2��Zw�Y�	�ʓ��Uj`V�kgTM�Wؤ�b�� y�֮�M�X[��u܅PG����wR��V��G�d���(Юr�
���lYT�8:�``�0q���2?��?|�	���'�	<���� �N��"vEέ���{�@������3�S��¿�@X��ws#%(���icY����^||�߃��+T;��j�yr,�f�_`������ײ��]rF���6����lkM�9�~��jgTO��]�����#�u�;��Q
��g�>A����{��.n���zĮƼl��~
�<3�]£���0���C�j9��H�"�Ji�.����x`a�*�W��S�	 �UZ�UXL����3�>��_;6Olib�u��La1Ӫ�»�ʹ�T
� ?�[�{4�����!� 6ŏ-~�1�.nV<�fuV��pg��L}!0֨4j���!Ipbxb�2���t����
:�$W�3��1I<Sh}�i��=h��B]�r�lTǛMN.����d��
�HƁ���<�`�Q�K�����(mL�f׼���$�y�D�~��4�%n�l���&;(ۑ�ÅA{�F_�l��~f2*�-��7���E_���i��X��dT�������<p�kdө�j� eZ��K�}���\�)dSn�ln�^�,�(v^՞غ=e��3�f�����o֐���*�o�<Ӌ�^(F,L�\
��(o�b�7�q�p�a��-��]��K���D�R�Ci>�6��N�<>�\��J,�o3���
u����2v^��"2
��t�C�'�[\��i��o-��% ^���f͌s�y}�S�m�AB�/́�����wJu��7��QlF7�S�"J��ǭ}}���X})�i�-��!y26.LAYu���	�8��W��Bt:������9h�e��Z�/98M�*���=�r2�
���5��[�JN+K�-��^�X"�!��� �ξ�i�wrP9�C�'��v$��[_��u}X�c&�.2E	4�w��e���i7X�|&$���7��~Ak��r$w�yǦ�R�LՒ�=Ш���jk��/G@6���"\�;#eo��apܰ���_h�8 �}���d܅T�hGυ/s�G����J� �t�g3^�!ݲR-�zO�JP���V��5�:T�+i}��v�'�.���\�_Q���w���nx�c��"i�7�C�����HY<s�z�lK�C]K��ݔ��܉���!{\�<3���æߏ�|\f�=UU�����b+�7��"Ά���3��^����1U.�p`�/�]ى����_-YK�̫�W~.#�M�dp��$��x��u�^�R��J}����@ӍEh�=��)맭����U�.��G�O�Q_��}}.��������x�:���7����n!�o��X�vP���D�xu)�>{f��C�F�p*�a��[_Nl�>.���������#x��`+O�i�)8k�ifL@Λ܍��U��%R_<��+O^g�����YC	G��������"^�C:D���fO2�Zݩ����
��}�h��?=P$�����:Ȏǃ��Co�C���X!�¸+��?����T���w�Rb�2��P��iw��vVDv�~�$��iN��l���9��.�p���H�Ҁ�!N����Z���g�v᩼9�[��>��|:���4�,������ӵ �B�N?�3f�Oܜ-Ա����0����tc�A��X[P�����*J���V�gpH2ES#�{G�w�vw�7�kQ�� r�F��|0��2��T�/x80�����6[�[x.�zVmm�t`�t���G`��cʶq��q����	y������"��%�m�d��&���F�f䨓rLǴ�k� �lB��a��أŞ�Br�K*�x\,>��G��2�ZY���S��~�m�3A�8;��ǵ�PbnE���B�F�'4��p����� ���ב��3�̟��'��6�v�c�F�l��0*�ߙx��F$bS�ӄ��҆��c&�Z����-�M�RY�ݚ�=>,!�髙�:of��|(�ߚ���~��E�}��l�
Y zɓGu-9��!��4MA�	�<A�-⽼�a�ʈA����X,�.'��e�^i*��cTQi�����	��Hs�Fe�iz?�^FeW����jF8�Py�ZEP,��~N�Mf*�i�\������	�����Z���vB:s�*f�z*�'��9xԤY9o�s��{�4E����~�FV��]p]Ѣ�Tі
=Uz֎�z%cW:�8՛$vI8P��m�q~��wF�|��"B�rvKP߂Y�<1�q`w	��z�3-��g;>kI�����5�.M�I�M���xٍoW�Q/����V{�_ �Ҁ`��5c">�ql�؆+�o��r^�q���[�!��T�6|��S^�e@G7zZ���+��>QsT&�μ���
��L����U	�r]��3��t�T=�B�m�:1�g(��V��me���m�-\�\V�(֝�ڑ簉	��cG��I�춪�!���5�Os:�ɚ/H����<.F��ZF�������5O�r_*ѹ5|&�%V���T]�(���SE,�+ٽ؋��[�,t��aL�'�1��o�f�Y�&���t�x��J0�Ҵ�b�}y�BڢrM,D�B�c�2���+��7XO�[b��%{�a����*#H����,�5C=��qUxJ�4y)��r�i��5��0���6�t�@�� V {���R�z�W�tH�s��T9��H���:\(K/c��TNv���=���Te�����[c{y����9:��S��<��绳�{%����.�<���;������"��e3Z6M����-��z�#�c1K�k�	�%���_�*�N�J��f/���Q�ة���S�7�8PI�����,���[����Dt���܉zi�VVa����y�8pb��j����@%7;o|/&c��	��	���&��)�׼�˂�I�`<‛G�S���v�=�j�3i����-�\��?E��7�Oq?�d!w2YT� ��#֕�m����)ю;}u��9�.}�^{���^��'��w l
^^?��vi��}I�S���r<jJ�̇I���BrW*S<6X��;[��ԍ0k�a����K�a�e#X�{�@U^��YC�ضF���iu)6���jI ����,�x�@=Co�)���y�a������mo*r]+#?E�����<���f�k����$���g���"M3�	�-�8�����NMmX�a��H"��{��J.�Vܙ���B\���=|4ѕ�T�*ت�����	��YI��Lfۅzس�m��ԪL�tЕV�ѫ�wM0�_�`O�!�Oa�]���څ[��χz���(QD��<��ڔ�,�#-�E���0��Z�N�)�XU����<U�]��AQ����M���O�@F�'c�W�/�L8x1�҇7Ϊn����ѐb�co��^8�6q�F1��8�y��x�qR��א�I�j�8�6V� ' E�YsK�tB��aNl~��_�oyT�n�f�/�G���gG}�e1b,�1j�&V��I�c�A�[rZ�5I�g�۰0�������f�����^���?�*N��|���U4�p�4�T��J!�}���kmJ��"�&�m��U��ਖ���V'�Vh|H_�Q���s���� ��՟�{[�.
t��1R���Ds����`Y"��	rn4��5�zbQf@�+��V�OI,�)�bI49VOK���٤��H9) �
s"��p�n2X��,B�VrJ �X �v=��)<ӫ`qF��t�<��%7�ܭ9x��@����Z{���w-(l2��<`Æ�G��C�c�sT��.�E���G�0Q�&�U��:��}V@_ �o��W��S\
�g=}�2	�0כuܬZ6��VMk�K�|ʖ`O��=zie�ٔc憟�/��19a�_e���s�4�׎aTRm�n~��<�[m��n��Әt�����g�O��E��!���[�cM��.99
��T��N��;B�����i�Ə/�4�EWy[Z\�(f��p���H�E@��>�Js����E�$�13���L|���"�
H ���\�B�	�[`0+%��Нԭ���bH��
�jGI�9Pnƛ�3A���:8�ڬ�1X���#�||eld�@��e\�3��]�l�.�#�_�i�0� ���&��9�HU�b?�AF<�U#��dE�")D5a9Z1{�T*޵\�sQa�tK	�|T��̌�E>�
�sq(0}�c��\��M��`�Կ�u�(W3��H�x�o����[���?�}ۖ��O=A�R��Nr���2P�����C��>_�uO1�!��t��/� j�)75\���R�˖A���e���f"R��f�(?R7κ�Yt���6&�h�]�?��Mli�姙�SܬG�ТKxA����x�j 2G=ˉ#�&mnY�|�����ϊ�u��F���Ga�Qˢ��.�~�1oG�ܓ���$�By3�_K����۳1$7�0�.��b�^�A6�by�8sG���i�u�S��h��̷���>�_2���8���:�����-�W���/h�k���,R�hB�e��X���������K�	��r�w���U�mBwep�˾�J����~Um3���:���Z��yr@�eh�%Ks�֥IF{z�ˀJ]4�g{����E���9�k#ϙ���N���߯[U�a�G>
�b�1��V,��rH���N�3tG�_��h����0Y�S����͌��{?_J8�+p3�n(P���}�R��NWz�~��u�ws�r����x@�Yq��2���L�<a�X���њ�S�2N�o������΍f~M\��IJnG��k����+n�%Gx,!�
2�'�@��'D���C��eW�B�{�P-��x�3"����KG)o*4P?��9�� z/�J��ʡv��{��s�0�H�}Hk�"��+�Z�uM�@Fv���g6#�2�/r����W��\+t��7��o�BO�O��<�	C��� ��^K�G�|�H0������n�B�/0�O�:�xT��c��4����>C�����ȳ��'��M����	`E�p�e�4N���1��\��%��"�7e��B��r��d��gI��`/�9XX]<�����'�$ݫ���J����OGB��ހ���;1jQ0����L�l\���Z�k��+/6�^�k�_죇��N<���H�B�J3oL�ZT�M����f��fBM�K8
J��Xصؕ�n���J�Ȫ4{�(ZYd�0�D a���Q�n�j�<����}8[�,��H�Cr�β�9�Lu�^����ȍ~��B��1��S�������O�ãϓp�˔<V�5Rk���m˃α_�S�pgû�W�$[! Z�v-.�M�I��8�N��|��gN?��52���Km����s
2<�E��(�]S?%���!k��G���:�ۇ��چ��ht������a�າnA�b&�4K���OO�[��J23V�%�ֹ=E֒������S:���a;	�0�t}�w�WW�/�k�Q�ť����6*J�]�s��� c��������b��,S�pS��Ϸthm�V�:�ry�8P�����cy�?9Xoc{&η�J�A$��&fp�"�n�O%M�w<�Xp1��q����hq fZ:8����>	s����Ԟ����y�2��P�0 ���ٸ���%]��HK��<�V�:�>���w[2X��W4����|)$}�����\j�k��Z��J��+ӎ	a��>Q�_���ë��c�{��	t#֢7/)f��U,��A�Kk���w(��:C�l���V3�����9����dW�	R$�aR²\Z��1X�D�_�u4P)�~s*�m	F�u/+Q\g:���y:�z"G���ě�����.�Π\���p�4��� ���C�g��<uv��ؒO����xE��P�X���ݮq�ឡ|���\&�f:�[)N,M��ߚ���G���**e{V�5lF�ZɈPo���*�`���U�5�W�֝?	Eݴ�Z��G�}�s����l��(�m��P���D��,���b��>��v0p�JP�ߙkr�{��l P���U���T��JA�(�<�*�@�Ҙ���cITAdr�'�J�t���Z�)�I-�?���!`�AG	��	�dՖw�mK�߅�������?�^������$0r�,�e&����9Ye{"b���Ӣ ~��b�o�[��N�њ�6�?@�"Y��	��>t��:�\W�=�a���m.�h���g,kMk�8� �j�E�
Q�	LU,�s��v���
D��ٜ�幯Z����Z���� &Ccvr�Nd����W�_+�����%9����p.*'&�J�]P/I1 S;I�5������`Y����HV��
:��W�A��ru#�8�;R'1�Eȇ �1aQ���	x��8B��8̢$.�+�)%]���p�/����ݾ+�`/�'� �9�"c�=�`rghs6�h0d��>#��O}�f�_�1u����6��k���GM>�P�쌭�5���m�f�g~ �+����X������.U�-�L{X���4F�ӎ�.���ީ=�@BQ��R�>��͟_���f\�����"._U ��gC���L����-7���T�C�щ
��[� 	�7DM,9�#a�q�m�p���4�r����A��w��D\�;c���W�2��Hϖ������������R�Lz�V�����{�{G���<>��&�8�Y.����u0���Rrc�HWxͥ(Sj�L�Fp4�EF>{��?D�ya�P �%W�h��մu��E��9$�n��_���:���$,���uya��-xNc���+��z�@����z�[���6!"�x~��*B[ƨ���y� �Ҋ�jQ�ė' ��3�.�@�����EKϽ�GO�3��S�M�p�TO-�����GzKɼB7в�r��$�òA� �j�����dX���=��7�iйS�M"X��Z������ޤ�,�h��+$Z�Ze�0�Y�4q2hh���K��;M-g_�,�%���<>�����cԓ�=/bK�ͺ���ji[����?�5�族6��Zd�|��3�H���� J�院8er�K&��7�Q{{�LRE��2�������O�zNڙ.1���`MȶsS�&��E��چCJux+���<d�Rx�W��f(,M<��"��|��#nܷ�R��l����F��Tt�՘����h��%b� �<�n"o�"c&2��w�<ȳ{T&��Tޞ���%$��:. ��\�eևa��'*�D1
�EDs1�*.��B�6��a��y���D_O������q^1S��5�<�8���+ !�绐m�~��������v���:�zM"#�]���ʞ_u� S\���#��F�p�z�����2"������ B�;~��[�0q/�d��>˳�+�Bq8�I?~w����-}sO	-�/FR
�lA�Qb�y�Ex�FA�hڄ��?t�g�O��P`��-��p�)�@�(�ih�@���:��H}���lc��	�L��d*S���2V�J�uJ��{rsx?�Z����/�\���M��OJoy�(F�݊���h4G::W��f%|�*=猈�[��%y�|Gq�i�U/�4�X�ƚ�p�o�yA���o
v�|[d�'�O��+�(КJg����Ś\���E��-SlI,{��E����G�Ξ�a��UF�v�}s��b�����AG�6��)����`�������T����`*�<���TLȷa�����qf%++I�>v�i���7}]5�.>hJ%@��� ��^�l��+i\yR�֚ghgYF��|?=&~*�����jR�J�f���"^��]X��$�c}��r�#�E����	�Q�\�J���0.���%�RX�����s�Be��ݺa􅷰��Jc�L�^@�wJV�jd����t'��}IQ�w�Jq��X{|XZ_�?��l�_B����I3e"��a�{���Tro�L{5��������b<�%#I���^��+��������αcZn����m��Ph��Mv���7�hC�����ɔ��M*k�:0�>�ZS�<�WHoV��b����ۯ�P���S�l���a�ݒ�✧��6U3�
b ]���ha<!�"��� 
I��W	\߷���u���2�)���Yv���>��H���ݹ��#�7�Kݖ���W�f��`\t�ȑL���:�����	���R�M��Mpqg�q�@'�������.C�/N$KZ~i�+O�U�<?̢y��@�(X�8M�����sܲ�����j�$~ɤ[�{0�=�r�􁨫�ol7Z��o���9wz$����#i�����N ���ٰiLO��V�2ɤd��H��v~���x����CY1
��ڼ%�I��C�+�;6Ў��=��teoc�`�y*��=@��(f$(F���á�w��E��q�T��q���FŸ�.��s��Xcdr����Y6�M�0���cb(�]����������������������:΢�Aɝ�p���~��|�C;������R�iH��rv�q��|.��(��M-13��L�$>1z~;��7=U{Gb��1뿷kS��ٰW��.$ؕw��{\[_����]sq"�d=;l��(�Ne��M�<$�`n>��=����q��u;.��!.}�**V-����h@�R*�F �����L���b=V�:8/{k�mn.N�}�c?@�c�9Dz7�{�o3��I��>���aܔT?t �,jU�=@����J��V�<EU�>�>`�h��G�4yk�b�u�϶}��-ٴ\ %s��Rݳ��>�9����}hߵx�廢H�AC�	�x��G,	���԰}��e&Za�m�m����M�ѲQ#���2��R��wD�B�͉�W�e8:OӇT�r
�	j;f*���:�$�7a��Y��8�	��J�Z�n*q>���n���r`"�䊞�}�&p�Yv��ڣ�}�e�;�8[�jUʟ鳵��ƗO��O?���/5S{ڃ�|^Y�E�|��?V��rFJ ��d������%r���{Ѵ��n�C;�g��P{���/ŵ�zܲ�5E��=��tmђb���W�x������ᔃO��6)�p?7R���S&t���g���C|dN:��(~u���t�i'�4���̉�K���L8#��ftc�7:BUT�&~䄽8-jY?�<]ݩ�<��tE�!�B}*b�����c�����:�2!��F��){��S:�q�9¸r��zB�H����,�|=묐�q�|z�����qہ{1�l��*�؟Lc����F�j��\��~}\^��xm�?lɒ�/O���1�8b�c0<�.`��ܿG)�g�*�[������"a�K��c�dµ	���;֥�R�VkG�yf#��΋MV6k��v 2�ci��:x����DV��E�f�|mIa�Z0Y��^�j��D�ʓɋ �8��J����ì�4"k�k��.X!�AM�Ш��;�$J�H�!^c�ǫ-c�i�K�{m���^�*'8����~���Y��HKW��a�Yl�g�(��siP4���I��'�Ք
y�N/]#�-ng�<��u�%!�}\7W��>ܻ���C��K��_2�v䐍l"k��C�N@�s��i!�C_�zLɠ���@� ���t=QZ�.�������X�ܭ��a��������ô��.�R�a }U�*J���$[�T��@\���݇+�$� �\�*$�������eph�f{��3�T&O�
޼7�7:��@�*	�Ry�h�<߯��22�'��"t���GϪ�aZ�.L��t�����b�6�ܷ�`e:�e�^9%�dՕ���?���xb�r�KB�:t��0x�|G��!;���2��gIQ���v�y莲��$р� ���㎵�KE$%K w6,����Mh�xV�uY�^�x�eL�Y6��C�U��v Z�.����^D�"]%G���#k"h��b�5��,�����&�4�'S4B�w�vsL)^bL���.z^;�u�N�ٍ��O@���$g$z(fuͻ�}��g��<��XY�z��}�,+%�^*��R�Q�����x���L�ιA��C{����9XE�}���%�Hfy�'�g�LS	W�}+�����9�T�w}�h�� �HXu��4��,<����s��]��u���@1����������c��B�Z�Üс����0*n��@it��p���$�֚��ƺ݋c�ֈ����bl��i�Ȗ�C8D�G#J��	K�4��>Ĳ �T�e�Uc��z����7�i�؈�6����뛩[e�s���i7�h�t[�V
}TPwڄ��-_F�.�礫#��$%� �8̆�
5~ Ro��������������ӂ�ąʠx�P����k3<0V7&�l 
�8�����c͗�������ک����V�O�v�X0��CCh�(���q��-\^�S2���?�<�I�V��G�@䄦��do�]�T!bb�S/�/-q�k=��N�D��7N]}a�F�Ks!�N>�R�w�MOپ����%�&d��G�2�5�ES�F&^`���v'�6���1��/{�Tώ�w��$KM]Ձ��7|�}H�bԋ��A�����ix�uD�5��1N�m �%���bA0B8���\��6��r9�M�*y�#��'�<l��t������:��jG���Q��A�r�S���k��%R��!6���(Ӛi� ^�{��⿷��#�#�u#�Ĥ��R4��(#!��~@Vo�zv�/�u�����m�B����5W�~O�E'ᐯ���YY}PU@nRT̽V3Q��幎����j��3l���ړ%���u=�'���k�e��﬘��6�rXB�TlI3V��M���\38�5�M��ج��.��*(T�D�^?��ȉ�+����"A�@�� ]�YE�/l9$R�+����p�x:H�V��+�br��aH��bN��+>dDN-)�$F��ͣ^�_4�\��l6�kHgTC�u'��
v��d��E�'�;�.7�����r�����7�x� �35^�Xn��΢�͙��'����.I�����D�$.��K(84Q�$3AfX�t�� ����+��M�p?�u@}C���ڀl��Ti���pt5aq��Ӯ�a�^�,�Z���93�Pl���.� ���f�@|ɛk',�	���zwσ�3Ƽဈ`���&��MZ����;�UB��S� �7�%	6���Z��+�C�Ӻ?%f>Ik|ƅW���I�����*��S���,+c�@�Ѭ��yS��5�,�M��e�B\�X�n��:�x���t��9h.�x�hP{���qf����N}�M�J�(b�uE8@bΖ�'\�/��\�A�߱��7��)8�H�e��P�:c	.;_�U�^��D�����uꅧ;����_�A9���N4��`*g�~Im�X���ݹ*���U��*<�㖝p�hX�g����q���M���#G�L"�?�5��2�8;1rX�+�pN����BN�����ys_�=��]�#+eA��c�\��݂�����c�e�%7��0����Ig��@�$�FK���C�aI%�i�fR�ŵ�6��9��i���p��prU��Ka�8�GP�QI�5V�y����)��
� _>��[�nŌ9��s%i� ����hY�tR���h}� �#|O!3?���cNw	�����:�;�+]�`3��@�S����Ȼ���/\bǼ��Y��(��>�|�i�n&=0�5dg�h���Z�n�庎 ��Mq�\��u$�b�T��G���G�~�xx��}�Թ��n�4\��뉽�x � A��nor����0f���FE&��]NO�\g��+�v+�fGnV��j�ʾc0�`��
�}�z~�oR1���pFu��qݏ�:�I�r�pr�L��~� �%�16fYv�5¹�ܳC��w�f�`Kv�4$j��o܋��*
�N�����Ac��L�ƥ]G鳖�7�.�_���G�\��d����Yt�w��f_G�d��5�h}���׀!�ѝ�j�g�xZl?U��iZk7NS�� �>��z��IF8�ӿ
 �k{\���@O��;�bR,�I�8�9\�(��9 C�5�s���Q�u`Z��S�x,TdA���t���&\2*��{"�K-q+�*ϛ�x*���P��p�N)�L�SP�ҿ`I�au5� �� Ay����mV-Y#�����p��R�7�AP������쮃J�/�`F��\���gV�"7��8,P ��)��M���F��-:4��^B �&1�6���L�<ˋ�������#��< %����Cɬ$�� �'�4YbdW��j W#�lTmg<����VM��rT�C�H1���B��n��R�"�D�W�ʂ�(��M5��_/� 7�	��.ܳ�6(�!I�o�$Q���kk�X5��(��b+ X�귏��D礋
@��T���2����@H�-�WlT��-�n@�b[�О"Z�7�<�b����w띉����a��Ru��?�l^�4��Sk;� W��z!nx$�G
^�� �l�>o:�V�/�=�+�9���(:�KyN�*�{#��sn"���B50��Z�p�]}��jX�MT>m	�a�3`�%�MF�GDi����n���e�ݟ�k�2��U+�5;��bΕ�`�,L����;t!]B>v]�����e�zǫ�*m��"��՜��Bk���cRx�]�q�a�5s���"I�V4�5��e�����Nv�.Pb��渄�ˣEE���a�C7�cnV.p���i�N<�:J�E�d���Mb����U�;����A��h�Mo�gp��mm�8���YB�M�����Ȧ��e��qν��|��<­o� �8)��V���W>�T���7��Qb��o�Q�{�G�)�.ptm@�)�#�fI��)p�L��Ƣ����z�D	š�����y7 �@�jҙ?0������sBwwWp�] @�Ҁ�r���&����;�N�	Ǘ3/��3}�
<�_89�;	�?EY�G���v�[7���B�'���ތ��f1?*#��0U�]����_�F(N��wӡtUn�(�M�[��p����U؁��:Eg����}����j���;tg8o���(�)�̛��>�d���x������\	7v{a�b�qZf��1��0Tih�ߺ?�zrhT-�PK�C�ꊻZHF�q��o������nhy֟��z��Ħ�Xӱ7R� �]���E�N�g����BM����,3Q�նj@� �^י��05v9�%�(�k���
y����[t[�jS���(̓��B=���6�O�#�g��j��~և�q$8Iї"��3�%�\pVr���k)�@\G���ە�מhc ~x]���1�ʴ���y��5�6�u	XD>�h�	�Z���Dۚa������,E�(�8�����[B�&[�S�A�م�iy��,�3X����ܹ̈́�p���h�P�Q1Dީ�zY��5�h�iW�e�y�B�Ip�S�Bp[_1PV��&��!��,A���7]6H�������ґ��yFx3fi�Q�nN�Ѓ%E�4��H��=�>��D��z
�Uw�n1�ؠƭ;��:���/yV��: w�+Y�� -
�F�Fu�5�����()i1?��$× $D��d�E�ӈ��kj���6�(�;s$J��K�2#���V�����j���35I�P ���EUk��'MK�,��Q�&9>/{#�R`��^3��J��2�10��|#�<$� ~��5K���?/�Qɂ��ረ�ʎA�\�9/%�˯H6�Q���i�W�fˊ��>Y���/�EY�bRp% (@�&Y�[�Z�� =x3%���,�</7r�b�J�:�u�yZ��˅����xJ^�B�}�_鼔�̎K�&�Q0���&�N�cШ�|�r�mS�y#뮭I�g�Vp�7�s4��M�l�S��P����U�Vm!�%z����V�Cx������ p�XVHW/'v�F���1;�[�cm��KF[�x�r������aM��.���<�t����A�ٙ���WH0!�\�/6��%]�G�?<������R�𶮳��V����8�Y��V�����kL��dB܇X�3'�vyu���5��S�l�bx��f��|�u�2=뚵�U)��AX�Y���.�{�vɔD�$f^�_tG|��y�z�Bȩ��lsN�
�k���C�cH�~7)X�j�$�~�'���?�t֪��XT�d�h}^���2	R�A�^٭OG�n#O��/�Lm����MUs ��a�vm�G�|+�Ma��̐�vښ�m'q˷�I�F ��r.���^�F��Li�d�Ou�7 �<7 O�5%R�O�ǻ��w�| lp�\�τ��Hmu[m�>���/E)f�E�j��Rdg��0�.\�5A_,K1���4*��e�F��	��S��D^��Zdk��)�W�MϢ\UC��F����u�׿�8>�fWj1�*(��o�9�p���G�
�9%-R��	jEO�i��H:�݉`�LϪ\���m������w�Wqa�޺pg�7=���/���\#X���l3M��]����Q0x���=��o�J�YW�{�/�؅�~j+��Ǎ�=�%��ׅk1���m��^?����K�\L�7���Gʛ��\V1f����Qѧ2Nh6����xëmfl���I�JAߤ��PX��߲��Bo��@*�hH���e�*!���6M�W��^� �ɺ7��[47�ޱXhi$�އ%v�~��|( K�9�W*l��7~�I��9��t���	�����t�GS����-蹓����PyiFg~�b���"�))f0��j$9�LE��DD�����ӌ�/�,k9R_M�+ib�u�.9�l_*d�_Z�}�Y�����|�s������OD����o��{�H�`����yQ�"�R�p�Yڂȭt+�:'%݆���,KP#���~t1�_<t_�D���ZR��%� g���Lh�҄o�/H��1����1��RL���A%����Tn;��[�'��}�h�����	g�m��!�xMr�q�W=�/������ll_����EѾ�J����� �N�������!j���3gfH����l'�I�* ����%��9�R��r�s@�� w�ՙ*��LN`شm��u�Yq��=r+
�.V�l�j>���.P���?�cz�P�:��7&p͂����ֿt��{���R�V�3;�+
`�
�|U��%���hz\Ti�]�R��@����mޔ�b@�S�O�Rz!�~�\�fHff�]6��7d����wUHpQ9#RH|�K @�܎��\E�|�<i �iv�781�pGJ���||xx-�,^^O�m��x�Pt�)�(��	V,04�M��c���{Fq�[�0��#�O�9������V��m� ��9� k��h�eԶ<�0�q�m73���{԰_h$5��:�f�8Q�mF���V�5���ɛ�A�Y�vi��^I�/��'K�Q�z$��1-�3e4~�ku]7��'\� ��~k֍1�:[�~1Y�x1"χ;�Ss����7o.O���'��,�G?]L	�N���\��>��Z-�yka3��i�o�L���-'�yx���������Tl���{��n%��:ȣ�4'*n��X����,k�M#3�>�N��L�\�Lfz��<]�� `@�:1^r��[5���װD��9%�i<�iC���yd��
]K8����1S!-v|�!Ը	7�--ݸ�g&K��QO�@��xQ`�w�]4���&;���������m�+�JZ������1\9�ٖ���@v�lA���r�@�²!��&d��
��@�ɨ� ��|��3Fv�r1���~ar'����:B�lN�k����Kw?S��'��`F��M�n?z�^�qL=��0�u�ўy�NkQ�b7��s�,��&o�Jp��6����\���q�J7�/�KA��.��u�#u���UT���3���<����r�>U'����s������3��p��Ñ��& Y/�6��&4����\Fн_u�f����#�ݑ�1�a�7u���'�c��}���]h|�[Ĭ��+�*|�7��$���xp��du�
rR}�֙�_k[d�4�u����� MP"�^襠�����&�P��v<��B�K�q��QW�qj�|�2|�c$\�e���D&2�H.��@r� 3E�>T����N_"�=������d���T��,�Bj���>15}�ۣ&���6�V�����j&��<I&��k��Ň��3eD�G�����.�n�9������oU���+�44��Iܩ�9�8ǁҶ���-���~)elx��&'���12�R}��Lc]��kEA�j�L6fEŻ�������h���o��&H�';
�1͙w��e�$#ڕ�Վs0U�t��:ЋrBP���Vwj���	\�/i�yzM]�1�F�\(?�+�4
��3����1o[�����3�
�w�e�)���2�Wsi�d��/�o�9�Q��X���M/�/9�c*�H:֎�,��oMڎ(3����(��9�K�a���C[�ʫ�({A�`�P���Yn(�s�sgg_h�~�]�[u�����O>l{f������u�ǔ�=gR��w�ھ�c�s�y,wkPu6�[��~��'��P�>��7�CKC���2�>/|�CU��n������\-s�Z��c��3��`|_,vUX�a8 �p#��qp�n��!������C�������6�db��>E0���j�`2y�̋ɲ����W��{n.QG�B�k?}p0���� �p�~�J���ؓn����6+7xg���3t^�1��r��,�l'[3!6x�~��5�*c�J �V�OG�4I��#� Fs#|-);���w.D.����^��&�I�*�D��09#�Z�>Aۧ�Ќq#�����`�b�������fӗ�G��v�G���/ͫ��Z��܅������jq������ ��$8��Vgs�,�hR,�k�1`����^�gԆg��T��J��h�>X���!*�|~���x�ti��q�S�]�ӟ������^���q-X�0;�ܖ~b�7	80�΄E���ϓq���v֞�E̡Y�`�OEYo��VH�F�ӏ��dC,�pߡ
׌�˷�B;�׹M�YS��=w���|�-iL�v��.�.Ƙ>��z���-
�5���7jEx��߁�	�ok�Ľ�ɟ�xɬ�{��Ղ��y�@ř�*5e�9��|����o���(l����r8Ҋ����T\v�E�g�	��&�@��BF��5
��B���T���b�oQ0��h��?;faG�z�����>��_�&����YJ�%�͆��*i��W��Z\�^��/�����gLWf`���3����5Y�
�q��)�K�ʹ��XQ۷e)��*�³��w'F���'_3x4��}���6O#�0�ܐ?G�RnuR�@p��[�%cZ9+{�O�oI����c6×a{S3�`/�\?�#b��x;��Ź�eP�3*�������L�E��`��$������?㬴���~�^�ݎ��*�U�4J$C���N�tLY�۹�ʦNIe���7�����Ɛ��&d��1;����e��)��ui��g�mMC��;��*��ղ��u����[1������#rEU$,��Wn0>O�;{�.;k7&�����;L�!�p =�-�����(��p{�w)�p-9l��k$Xf[������)�*��5c��Bz(��w0�i;�������J
��&�[7Z���jH�Z�'��҆�T��n��|�Io��&������)Q:��v��C ��Hg=q����~��ǰϲ��,�uH�lr��``�7R������Z��y�P�A��T����Q����-Ŕ�{�Sӏ���f��OFc�W�R��`��p���l
�\ֻ�N��7�o���4Tz.PUI����sQ:`ִ̚���)B�qP�+�Ue�J�0�*H`��1`���-��+k���I2�{+�,�2ߔ@�����2L$�m��{�>�5��,dJ`v9v`�Qh+X��{8;���Ɉ���x���Ȕ�\����o!z���XQY�ۗ���jM�(�pK�X)���4v{=��KsE�ڋç����c�w��y��6�J.7�`U��ʒ����Rsy�@*��N&^�JT�4��[�q1	��#��O�O<Tƥ���=�Vy��[��� BK�8B����&=��޺� .tJ�*�q!��!�9� Ѐ[�^ՆnR̟�;O�0�N��*��k!��1��e@B��Ή3.��c�m4��A����X^	y��]l�%p��*�eKcNX��&� ������ꚗb"��4�3C�O�.��#���T,jsР�Yp��� ���|��GF�����������"L*'
��U�>���8��ޗ=�p!��B�qء��Z
3�d<~a���y\�����K�X�/ʷ]	��#G4�}�T�[�
�	)iĦA�W��,s#mG�&I��*�t�M"�ݤ�H�>~�$۷� BjzQˬ���H�q��������T�j�����G�q'����C�
)�D^�j���Z0��S�U2γD����?�����ڟG�h>��+~1b��4Qs%�>g�Ri���+���C�%J�<�jtN�^q� -�-05�u�1|�[jG�W��/�-�T5�0��}��3v���Ȁ,;%$�0�"�v��Eoxo�D�$���;����/��u���(�{�G�y{��˒S"�V'	�����d�4�R��in�� ��-B�I���@�z������eC� �+�@ȏ\�+�ycB� ׯ�v�Xq���g��M�Lj ��\eofDmP�Oԁ&���|I�\Y�xMm��ΰֈs]�e����U��
`�*�����b��a����ٱ��u*�}t����:S��<�1Y| �A��0�(� �����C���a�HgI�0�\�>�*C.ހr�ʹ��u��F�1Ϗ^D(��Gn����FR��܀᩹��qo'�1r�;V.��9gPF��Z�Xe�XӶ����sM�K��I��dJ��#���7���)l&�6*IC�F������Aص�;v�4(̵3�N dRو�뇥��.���	�)�wň����#�*�o�g�j��:g~G�\f.����7�߅��+�a��"	�q{�R�hn�E�q �d��h�Nt�����GETG
�g�P�nx�- uX��� �׹�Ϟ�vg���㎔�W?A,[+�#�7���yA:���)/�!��< H���"*=	�P�񓐑Ґ�o�G�.�
����E��83D���~+AZ��~�z���90�l)kM����b��w�U�6�zn=���P�E�,Ua�����,����4����(WK,B�g\�0���	�Z��`��MxU ��*��&�pZ�i��Ot'�vt�24��d�(�wA��|?+6�ό���!�錜OT���p���I%r�����!ԅY�p��H@
qcW��#����';���"�d w�*����ݻ�}K��9�X����8�|�溣�Lk� �@��g��p*
�h�w�A�����RǺD69��J��c���M�D<ؗ�`�n5b��h-mM_*����+R���\l���K7�����,��h��Ecϯ[��_��� �Br݇� &ȁC)�T�->�6�|x�������p-��&��ꀠ߾���xO[j�&�����w��4Vh��B��^�N��#���Wh��3�oN�}�!���	�j��'�6Cʴ�E��Q����ޣK\0���3�QH{Ҵ$�m�!q&\``�r��PLv|�&*�q�l^~��� �Ma���/���L϶-Kp�j�/d����0,}]"��s�"�ω���������tC�]��!�?�5_�J����ҵI�ϏV��?�k��Q+��b7p�Ȝ%��w��񰽡���o�Ʈ�E1s����`vuq!��������)a�|X_gW.+�)��QY����{��vi#�>�b�p��wͥ�����hD�p8g{�ˏ�l�ѥ�"-/%*2g��%�U���*���='/<�v�֭�����݌�蘨X%g��2�	����`�e) �o8&�wAw���� ��G>JZ��~(elS�2o�6���~l������{�q��"
}F�P7�#�RpԶ�SU5��:a�]{��\rP����y0�*ιR��&\=��%��}[�vCj5?�21�7��������+���B#yc�wѷ�-q0[�Y��`�;Ǣ͊�XUJc$��٬v���0u��R3:3J�b}����D��[)�O�W���_MtR�7�-��:nA��t�|���ؠ�`�g�
i���3v}Lk���uq�;��f�J
(Q�����;b7�A�:/��v�2��`�1�o4�=$��E�A����7�M������8��9�æo��@#X� �>�V�1sJ�w�*������:��v��l3pj������	D�x5_K4n��v8���������Z-�8{/+^��2��}yw.
�4<t«�u��$����n���I�{�H���������|��'�2�Zb��]/�S��=Hm�3��f]��d��
��S��1�r�?�2};-�ȏo�ZG��]�����hg�� :͇l��� �	gR5�H
ik�oǋ��Rט)�Fb��'���#���׫���-{N�Z����K�=YG2���+p��:䏰�Xܱ�|��c�Ql�Ah��������-?a,G3FW��.\�Z)P���);e5:̪������f'����Y91��0@�7�����y�U
R �^�!n� �W��M����-���mr�J�||�6ڏĵ��W��	�>�����Lơ�݄��E
0�����F��l��E�I��*�EG�NR��P�WIT�j ���$k��PE�|	��<Z�A��q>G8F�����׵-���/bb!��=�P౧�Z/SUR�a�_�th�h�\6� ��C(�����'�����W�&���-�����i������Z�D4Nr��N"T��6�D9�hy����\Mh\���ɯk��>����(�a�/��\��:�f4d�4m�0�,
W� ר��B�)>�R7X�}����Mb��	����&��%�l���=C	^1���%���q��hM�/!`����
!�@=|�U�C�z�0Bƚ���nJ_��.���݄�D���h���/Qc�+K�٣��>�9��W�g���쳥�	��Ў%<:g?�G�CS3;ƽM����E.����e ~��@17\����j��͵��5�.�h��Q�Ԝ�*l�a>�6��(�B5�DX�?ВG_������i�-�_��c`\���e��<�o)u�GL«P#��N�d�K��.١��1�y/�֩n�5S+a9��Ӣ�B;^6���L{a�Y3��´0�%2\���	l&��؍&�U1o/�yYR|s�c�ԏ�5�N��Wa��I�-�P#<�gv�#ay�����Z�bfr'o�(A���B7���NWt!&Hk�	�����Q����w��,`��2(V�g�/���U<�c`���37>/��\���-�KYv;/~��`��{���93��Ux�U��MUҋ1et%Ë��}7*������j^�V2O�~p(:�TR���X[KJ���ۄ�)��W�sA��f8�.��h��~-w�Ӕw;dH�f�����w�繖+��h��)}�ywuc2�:R�])�AV�Ո>�Y���qCPd�2�Rqkt0��=�u��L����*qoN�3M}���� ��`�p�Lv\ͳ�uƔ]Uٝ��ݳ��L��[	��1��9���{Xi�;a�HhR�vaOK^�^~�e�	~)�d(���$H%�~[��q��5�$�u��Y��_��&s�7�3��$r�������[u=P'y#��W6m5ٞ���4"'����k��<�獵�a�K�]��JU������}�'��(/s����f.&��J��]&��ƨ-�x@�փ֑Xx���U[N]<Az���
��ʄ��%�9� ��%��QKP�~��/�k��"�$ѫG�]�����l_$��) �wT~����aÀ�ĸ��%� �;����w�^髫eD\��Ú���ksD���Mgw[��N4lw.��p��k�0���7��^]�'r��Z��X�q����Y�Z�u]�2�������a�Ƌ�q�bj���yp���y0Mŵ��\1�Cg��_�������Q��g�]`M�-�w1DM+q�ss jbA�������'n�����˙�̖]lij��[b�(�vn�4��S��rŧ�uQt޻����Y�3�`��U��NH
��0��h�{B'^ksy]�}��=��v��x>�3G�=�RUk~��*���+�n&ї���ĕ0�E�K9_y�QHƽ���9yf�_w�jf�<=z##1������w1:�E�z�ջ�~s:O��zY��?�
�~�f��{�Z�XU�ATI0�tjYF�n7v���ʨ#C�=��LGTmy�o�Ͻ��W�	�>q�p��_^���ԥ��yK��4��O�\�z�R��¯�yA�(E�P���
�-� '�8C@e��1�W����Vc��ni�b��sb���B:�G-�f��7���q�o�s)c-!
���,7��Ŭ�f��F�)`�ʱ�ܪ>�yr�4�.1H��OK���I�d� Q��I�o��Sz�a�('&�9S�%���K�����LO�b�p��+��L�9w'ҏS������ ]��z�a�Fg=�w�݋6/��{JD�Ɲ%d9oyl-v_��8���X;>&�"�+X(\�	rUL�n����:ߔMD7�ym�)�F�D��WbV�8�Z'wo���x�ƕ��aLmg�-�Hi���8�����!Q��������2��֥(^2���o������Vfz���i �7'S��8#���Z��VL2UϗiY{L30��D���K��|/fd/�)�c�@��Y�SGh6fV��&à���~+�ɉ��Ғ�ZX�65t�
[��9�JV�r�y��|��ߩc�Lx��6=C��v��l�n�;�@̻�5 �3q��@W�;���4�
4ѿ3��d1�Z��5�qQL`����\�832阕�IbGjl��83�Tx���F�w���]��B�V�Bi�/{�#�l��y<��-��٩����b�Y� ���b�dŀЉ������0��`�3�,�7]L�̀J|��bZn��D'��x]���;E�d:���k�[�&2p�(��G�[�X�"o$k������y���o�TOas���ME���1/wa�;���,s�8�����	H�	����x���H������Ϗ���Ac�S�HXh	������X��\xB���jT���D{�{Jߣ�b^�P%����|�fV���A����h�����o%�ncX��Y ��CQ&*���I��pL�lO�q�l3�!�"�w�X�v��Ϸi1�ܙ���Di�7��A�3�{'�h�֜��!�8ONP��a���*��N~�ۆ;��'�R�II�9��_M,di�@vB�4穦��b菔J��V#x��E�|Y\c0�f�u�ۡ�b��L��0�6�ʺ@wx�L��������
Kt��=8��_p���ڿ������M5��X��{tN	�M�>a`q�r��N�6pc�ps�8�����H�S�)sҠ����*K$!��HDs�g�wF�A$M߿��J�n�N�1{���U�v��nF[� ��*tY�n���Ĝx$y�$�0ĝ�=��f����a��ik�Z�wE�Ā�&C�������*	]`�-�={�IB"�?��1fg��!`Pe���Hs���'n��;��'C����B��C�'aTD���&����{�}B�ǈo��w3v��1,�sh����Φw��nv!:�w�.exm��VR�m���f����ፌ�����('(��z0��m�<OF��!J�?̽ ��?�m������$2�4��J�D����U��8��"��W��WYM�SK�������0B�k���[����s�<?_�F�x�ɕ�(;�)�W�]�&��ӊ[�.���h_ ��CK�n�i̲�ӄ��8��/!\�j�	ml�U>���*��ɫ����M+]}���	�����Br_���mk��EƦ�EC�N�{�Y���=ʰv��c�bO��bg*��b�ž�  ��K*u��Y�$"̒�eF%�{0M�j���s�TY�Y���P����-Lkq{�ǰ]5��}���R\(D���MM�@vn'��-�Z���8W�?��)�4�P����������O��6���j�t���2�}�}�+^Z���B]�z���W�$�j[m��P���Sp�~Sk�swF�t?�Ԩ��x#N*|�ʲ���1O�U\LM%.�0H���НxO��7�����#��@%JzT�N|����q��DU�t��;��jW�L���;�1���و�<�aG;���i�C��3Y�)�����v�?����<.bՑ����\)6tP�o�TN�

��x|_��}F�;����Չ4�BOg|C�F�=��{b�4���d���9�/�*��fOҏ ������� �(�V=d����^�n?�vSL8��n����ض���a7>>t�G���1k����ý�so�_y�V��)$u�t#[�;��>��D��A9vWЂ���2��s����|(�џџ�d	��n�D��7����Q��%��=�rQ���f�rB$��(Azr��쩮~���I5�lE�������������c��\�lgeM�Q��NK}
ǳ���zD�g�#/ζ#0����MAd�T�8��?Ë�1'�j
9���U��w����F�-�>y�,ۢU,97��j|d)���C����zxP��F@2P�"T/Ӵ����|�����묈'�cf^`W�Y��r_�r��kQT>%u!=�嵱��1X�|����vRGr�Ei-��SG�a�y��'��IhY�����TN&�B��f�s{o4|v
�Z�g��X��N&��di�i��+hg���(�8�%�X����|#}�R�I�4G~�u��/�I�A+��|s#�#Sq\�w"�u�_��xqc�]4��J��+H�ѥ��c���	iѯ����.j�\�t+t�<�Se2�+�e�D��-�R\�L��;$,~��g��UM��`���ֺ_x`��kJA�7�m���b[�2��l��Mt Q��,�c�JP�)#θ�>NigakN=oZ�e�nJ�z�$�' G���n��4$��6���6�Ҳ5[��L�U�{vEV�j2�;����i�!RD��	��ԣq�3��j�=Qe��&MC:D�&�o��g�4��pt�n��:y�ޱ;�٫�z$]�p>����?�*\�D�G\>�s�������O3�z��HV3�
%��������6�"�Z��/m"����Ćx��(���s��7����xʶ1��Ơ��z�w�lԋ8!��eQ�d[Ь�Z�ā���b�a-�o[�`}�F�럖nQ�.��:����N����nY?V��!H���b�����,�mY��e��E/(�f���k[)U5��M˷����גI�PL��%���2��V��%{b���S�g�Um�խ-H(�@�V�V��+�\�nM���(z��ʢ��W��`�i�̢���
�`WpK����6�$�`也�*���&��F�*�rA��])�"]���>Òf���|�ʦWB���x���jӥ��S�[b��$����3i�
^ec\Fe���(� g��8DP\���#��_����Uz��i:��lT���GLܲ�5�����9����6Ί�Y�1*��౪�F���ڴR�&/F�:�Ҕ:xV��=�2��R���w7������8t=�N6ʵ�N�o�a�����`�ike���d�����v�^��t$S�D��_|��ƭ x�i؆�h��뮕�2����q
�n1~�CI�V���`3�M�;s.=�Qo���}U�b�@g�ttk��_�\U���C�/����R�{������P6��6���F��o�N"K�Q��:��� �� h�vW�#4�64zcfYڥY��~�z��+'HB�;)̟tf*Elh�wL/���(�Q*ŖB�!�"[�M��va1=�D�����tP��q�ʭ�R���F@�#��=�+�t�^��Wr�(��4��,+�J�2=�i+�wp�v�U"��"�U��i��Em~h�ָ��]��7�TXwk��Ln¬j�/����<�Y��F\����A��-�)w�:,�
���(�}��ZG�呡���ORӏ�����ŋΈ�"�m��-���}�[L�2�[}���w+dB���p�6B#��o�d��y��b�~�Z"9�~�X��(NBz��x-�Waޏs�����[�T��'e��^��2�/�5/i0�d3�	���):��izK3r�`�Hn0���wi���K(j
�i�j�<<�S�܁U�
���h��u�ڵ6µL>sV��n8��^���s�b�P}��@�f��i�z���u������%������>��9Ե��+���WU�Z�h�j�/쨭���&�L@��6ı /b�IC%0�ʅ��L)itn�D�F]��v�xx��JA�o\�ϽS��
��IYްIL/,�r���&�SG���˟�������?�٥71T뜪u's�[�A|ߢ�^��ֆ<q�6�O��L���uc�} �2ѓ� ϴ��~ב��'|�G�k�@<�ܷ>2��}��/04-�K�{`���&ǣ�|�+��F5��dཕ��_���gG�˿�LNY����U�عX1$CG��6 ���//�ec-W&g:y���](y�/U�Xw6�����=%��ʀ�Ϧ0�&q>"�[ ���s���Ru�ҧ���돷Ϯ��,>qx�C;>S|�H��72���N?$�M�ި�g	���Q{$J=��&�~�U)���@S ���ll?�`�c����:� \#4�5��L���C2��Ku��:E�>5��`�2�SUN�Z����H����?��s�jxGoh}B`��(�":1nk�xS���>lPv3;�JG���t(i<�lC��e$����zG���k�5��-iJ�4��<��X�Ө��aR|C(N:���& jj�b�A�$O�S��n��㲵�_	K� ���~5"���Y�NeO"����I�9L��zU�n%�I��������RN�BJ0;�z_Q�J��S5�_sa�>��������}#�!�ϼ��s�wX��u�J�A��_����#�������@��/l�x�g� P�0��Fq�3���
��:��)�l��<��Ha;��S�S�,s�[��}7 ��H�u������˺���.�-�\q:p=+��&���-����r ��Sr#��3�ܺ'rU�}� 6�+'�g�Evw��>��ґ�_���n�~0�<7�>h\E�)��&IO�$}�%u
 )"D�y�VX�)�?J��RӮk����"	u<���"{����Iun�x���d_�\����6� 溶�Y{b���>�1�>}Xw�>(e�*?�T��Wa�������P����M�0a͙�H#?(u�0N�d<<��G����c<�a���j�4+)S:d#Ft����}6J�xއI�C۩,��,J5���`�'6�����$�}�Ƃ��nQ�u�c��5�:�fQ.f��.L�	r�&-97�H{e�ĕ��=���IO����=.�!לrC��z���]�|j1��0@��Et��=��q:������{�Dql���n�Dz~0y�q��$6�����GF�D���vg���r�	�\X[��zG�sIF�q�p�Q).."+Ԝ4��m�y���̶�K$��kѴ,ݻ�@E]�'���[���=Ƥ٬�^�ݕV��P֚a>�Ε_y7;�i�,s�@�,A��6�y�_�������wK���kɹ��3�W�S�}	���Y�O@�V7��=�H(��Ma��G[yH��M��W&EuSh�m��1G<�Q�U��Sύ�>�����ǐsjX�[�BhuX�Qގ�b�xK�gwM������M��� n�
k-}(E��2PGqY�Z�l��-x|��ӥ�1��= !T�6�Fe��N_1)��ڋ�ys1�����u�!@�S�#�?O�zI���i(�8Hr��[�]�7`���a�/:���N95�\}��K@�G��u|�^��òa�>Ȃˤ�|�&�BZE	T�wK�(IX6>w�v��Ӕқ�b�IL����h*��N��&LWb�?��2x�'�ț�{��L���w�e?��[R~l5r�pDD��B��N�Η��R$P8����-���5(
�� 5�G�ا�>c�$ۇ�V}����+>� ��N��vӒt��5��>�I�02)�>���>ZFcצN����no{��c�*ƴ��f	������`�P� �t.h^�)�a. V7�y�N3�0�(�����Ë"���C	&�tcY[/�k�ŋ�8�KBHKB�m��أa0��;%<��ڟQ�R�U?7׬�pL��P��q��!ܢ��f������(60>|��~!S���u/}:���
 PD�O8��Tj�,]����=!E}7�~�І#5�7� 5�Ղ�jhdi��no>��L�ߣ��@E��V��Oo���պ��]��BP�jQַD8=I�y�y�����niĆڼ���j�7K��lC�-jT$3�W��Y�2�0_����j"��IZc��[���!u����V��8��
��4�\șYN܌���mD v*u(���Nv�>�����]T�칺�p:�]Y@��j�ӧ�oU-Z ������غ�����t���\�ש����^ ɖ͛q��9ԇua�
�Ƹ�D[��Y��/K6u�����)�2��-��Gޱ�D�¹> ��iKn0��Fcȿ�K|�Im�h=��}l�UR������y��k���,S.+ҕfC�A�Er�證Ȩh$~E|޴q�|����"�A������v�E�zq(�x�c�8�4���^f��\��.��z��*DЦ�����P�/x�����퍅Ψ(ԗ�~ݜ�v���l��"},p�A{�̙�x��YA�+�s9TZʮ����/���|��g8��;U��n��2���پ�G
竲��B�7��=c�n��O�0}`V�=�d������ ��D��#3K�a�-p��=|C6��'�oI$�ȯ�v�	?�� �2c�:�ύ��0�-�0$��>��＿E���f���? ��c�+��F `z9�F���|;����O����:��oŞXk�c^�ds 9��lKM	7;A�ڞ�<Q������Q�&� �,�Q*���({� }(�F����D&��k�����V�&�-�}fH,"�IV#�{���:����n&O����`/�s���J;��QK�#�(<̨���Ȅ�i�;�ʪ�b]h�EI'���/3��f���Rzgh-���⤦N�K�2��]�`mX��K�?Y��Ϥ_�ȇ������J�r��z^�{,�w���c���&�G��a���b�PsKsҴ�T#=��s��ᄥ��ly�1#�#��d�M�4}��}���
0E�N�1f�) m�<��/���9�*L�ޜ.���~� 2+QE�9J5��x�FJ���&OlF@W�O�''��H�������83~;����| tm�� h��N]AÃ��5UZ��P�7�B�����U+Z��WN�D#���\lniI��
0��2/{�ͮC=l7��My�0�j�`bDv-?m�����v�)��� uW����8gt��U����_�����P���N?�I;[,��?D\�˓3zL�yY�z��[�2�fe�1f���:r)�>a���N�<����������yߺd��fP��CO��#��TJ��EU�˶��֠c=�O5�}0o8W9觏f�Ѱ����y��r+��]]��`�ҖG�Y2���X�ߢ��*N5��G:�=͟U�1���oϬ�aL�;@LY��H�g� 	3?`��S�%�ë�k��-Nߵ��Yk��-���������>6�~��b��܋�O{)�/ʽvk1�[��s��p�_L�7&C�<���Uy��b��Wc�VK3�N�iW�Nb�d�}���9y�"{��*h�S%H��� J����[\!��ݣ�䦳ῡ=�t�����~+F�o�G��),�%���&�=�X��7��"�L�{��kHϯM�����v�BՅ�?
|�,�jG(�!A�t0�I���g����:ٰ�ݯ�yA��gK�����)�Lme�K�%�N�*�&�vd�l�}�#3���VI	Gg�Cn�|��\:�m.��{>o�����gaD��E?��_���n�4�dD"y�Zt�4j!�Ŋ�'�Ս�Q���%)B
�F#Ka�m��֧�*g�ǡ50�ro�Ѷ��̶hU52 �+6+H#�����Ts�|�g���{U<�q��_�����=��!�6��+����
���z���5`��!����-A���L�3K�(X�Ldˍ�'�γzy��:���Ǳ���`��)j�ݔl �G�]����iH5TEs���� ��
�w�m_�Y6��õ�(�ƃ�v�����L,A�ҳ4�p�#�D��5��`�Y#,���(�+�〪��X K�Tm��%�w��H�����A��I����'��L�BA���j�:^원��2�f?�"|�Q���Y�mO=%o�3m�6��m��� I�*��kc���pݭ��L$� hIv��z�q2|��N�K��AC�@)(0���h$}��.�����R��Z؁�u�F����9!���$�y���V����Nۯ�}�~=~�~��b�����2�@k޽�X�ڀ�l��#��^Әw�L�en����^l#�,!E�KKXcþ
H����Jrm��JWeߕ�͟�2*�(Ρ���q�Fؙ����q{�K#(dݨO�5�5h�������-7=��������B��g��ܷ����>}�h��(	��a1D���F���b��<3� ����Y.R�`����-F�d&�G�ESA2=v�xB�!ç��Y:�F�͋���M�����F�Ta
��~��(�Q���W��a'>r�O��b>��) ��_癹�j�Y�ĩ:��F���<��M�	�մ�mI<�*n�� �м�׻���1�H�j]XQS#gǯ�@'����ǩ<9 Ψ:��;�bL���n�U�]m| ����ȩ�G����(��	�MEBq�O�G��&��4� oMu����HԤ ����Z�_�3�}�.�7��l��C�X��Ћ�������bAf:���o�8�='��X|�}��ɶ��wH�r][- P��HA!&3V�T����0��z�y���UF�2;]�MI��(Fɏu$�g�]c�2�j�"�Xc%F���຦�5�����R��] L($�n��z��Ni�nO��2�⊓%̒\	k���k_�X�	��,��42cU��fq��T�T�WW/:��Je"$0�%���M0����M�#ov3�,����X�*�S�K?�I�'z��lm�׉�^k�A�sآCv��/X̔Uq34�NY���C=��/�#S��	k��M�<;�M�r�������:\
����Wq%sa�aLu�7�M���k=�.źUj�K��0[
7��ò_C���)��w���H��5�u�x�b�p�H��z�2��Ή8Yh�Z���&�G�7��&��'5���9����3�F��������N����F�y2�,*�� 3$v;R���K�6���]�]�����k��k	�TM�fty"�<tW���
l�6B��.-����vD-��)G�v�!���&��:zV\젔��ə��v��SZ�1�C��_��Z�~�XEr81�I�tzU��$2�l�)o�d�Тa#�Tf�Ѹo��E=�ښ�征�iW�	J׌ᓜ�-u��pa6#�|g�HE��L��}�Ans|Z00>���d�,��\�iS~b�>�X���vnv�7���?��LC^������b $��:)2p0��̃1�DT��	�J5׉u%14��eС���_�c6'�2ߙ�.�
����u�����T&\M�*s2~�>u���{'�eL�=;I�VL3BG�wT\����c�fE��\j%�ʉ$������8 qdf_�{Ё��y"3��l����Xs�D�mxD\z<8@/aH1����7(��X_�w���/����I�D俌>h������ݬ���c'�|�$x�$��$�$'�@ŗ��u���w�\-�_�������W��8�r�q�r9�
ϐ�3��C� ��� ��G�vB��4�W��W���'8��J�B�;٥5n��
K�Dp��]�#w��A�P[���X
�j�r�m��Z���es��|Dw�?G5�:Ѻ4�r᡹H8�n'���{�Z������U���W��;n��\��� �A�|��S�5�r���`[�l��4r�n_���g��.#j�/�n{B����}����@`�]�������E]�~cػ/�hw�����܆	cE98�>��8?m.�q��ĕ��d��V��Y�v6v+j?G3�y�	g�'�������!��!���F�`�&ޭ�4RUw~�-��m�8'�C�W;TQ/���V�}1�s��f�j�B�49�F�F���Ĭ��\	� ��K+9��=B�G�U��Mo���,�%Zhq�TCW����80z��v7Ўگ��K�e�qm�3�%�ESs_4�(�r �ԇ?b�A��;6�!z�IШ��b� Ʊ��
#�r##Q����3��ؙ#|_��=t�a��4� [�v�8T�n��2,��!��U"@#��ɏ�d�F_2P�~<B �F�E�\ ��㞃�t!H�aEP���8�C+F�msO�?���c���êS+���[Q�php���u1xF}g.�$�-��a*�Il�6x1�|x��^�V푻�7"�I�+О�(f	�V0tג��PB���Oi�c�0�kY��*�Y9%�G�����4iC��NVC���6Y���o|7�6�jB�Ug$��TU�4�!Q��F�K�T���*�$e#q��>��2RsYRdIk��C
�]���X  �'��.SD%�	�����H,<�,�|���ذ�>�[�A����Q���x�Y���� l��$x8:U����͉�ˣ��e.+3X�Aʾ}i�B��Oz+��ځk��(2��?�6_�W�(�]�v΅R,�#h�6�H��*�W���q�9�+��N��{���{����5�Y��GK��:���:��[�̏0	o��e�F��� �0�SBƅk�c1�
x�=5���hT{�ʑyP{��\��;3g$�yi�E�#��}�*�����	C�����OJzB�������0cU�2
U�[����8X�6
��F0�(NC[�\;9�ִ=��1 Tv�F�uo{ɤ�ϑ�B}K��On�y(��6�LL̪�̕�V�Y9�P�7�L ��׽9>U�˔&��F��]-0����</_\?�p�!e���,��}Ǔ*��e�9?,�B�_�4���yi����(��!�u
GT7��Lw�4��I+ k�^�ADLZ�o�BB���蒩@Kջ0=4O�R��Z�x��I���v0֋�f<�o^�4�r ǰ;�`a��j��AM����oͪ{A ��S�`^'q�.���#E!2�n@��F�#�a߆���	�ϔ����%*�|xD��G^̭�ދ� �N����^S�-���)�B��64�9S��>_��Z4Чz!Pw?ӹӎf��U2ގ<N.�1�x~.�Eo�����&���`-���bu��.����Y�f��XA�.��K��u  w�����8���������%�s� E���b�5��$���a�xpR&u|8&ٵ��4�������)��2L ź�ga%la�8��4��^q=���]n-�/�Ю�
 鷽J澦�,�?ζ�N3�@(2���"��-���5m9r�8��E��J�Ӗ���B�R&���Z�ۑ�bб��mv����m�'�h����Ǥ���4���.�]{8�7�ɾV��u��z�2��H�8J&�ݏ��#]A��JD�u�����IQ�~�o�x�/���Q�����g֪�����ZBH{��1�
��ìc�!��d�@#��Ɏ�r^�e��L�`����?��u����÷�!��{��"����N����?�h\���z�x�E2���۬�r��^���F�TM�kK�r7&�ȫS�C�����%�	��}�-�4�3�B*!�=_�o��9J�7篪_�e�%��-��q_T��e�Y��$�b
p��}��^A��5S���5#G�\u濝�X��n�-ݷ\��O��X:��^�	�ѝ�8A$����,2L�;�&e'�l	jd�|�Gӓ��\iqqs�*r�^_�1!U�����ƑG���v�kǗ5[R���=�S�@!c/��Q;�Y?I\�
�F�Hwx-L� A�`~(���~��{L͡e�3āǒ,���p�5�6�N}?5P_nb��e�uѽ.|�
,k�gu��DqķOQ0�<�-�����#����p|�l��A�W�լ�Ȏx9�I���#���7#~2-���d���"�&�X�|�V1�($7��S��e�$[}V�gԘ���\N�
0��,&P	�-[��p)^����
D{�/��n�9���H��(u�F�K �?��v���B�;� �r���?e��yk�M���%7���< ����x���,G��BIq��P� A� �tc��P��3�X�3���zUhK4�N�]Q�?2ZR���� 04���<�]�S��Oi*N���������������y���C��=�U�-����Q��59|��¹ǎ������1�!#�\�][�>���5��x�|�m���/n%��	�܉��!a�k�f�N�M�*ҏɰ\�.vˑ1���sf�	p�qyk<����P��ǎ���R5�loM�@�θ `��g��`��Q0o#-��g��Q+��q1l	m4��Y ��-}�yv���kiC���u��*Fwj�%�P���w�B5��M�>���o����X![Y(��` j���V�Hs�� �&*������6&��}�'OM��l����>G�I��	J!����ˮF��)}T���qny.�i0�v�󀏱l����r��˧�_р��Ҁ�����B0�]ˈ+yw���yR�Ʋ��Sf�J�o;��#�hf��������ҜWF�vx.7���g�I����GەH�����&.����G�b=<�T�Ǵ3�F�ȋ�Yb
������r�2OT��0C?&d�r�t�%�Sy�X�����46��WŋJ��:�+�;�٨�J^H7y����AW����tbs��O�`1����a�h�[�D�w��;y�h���s�Z����yR��Qv��V�J�Ʈm�� ��L�~��ڻ���2p,v���H&�wԢ ��|v?�3�7� j��5������g{\�`6_�4y��>����_���|��H @m�}��Q�ecƜ����b��Z\���� �&a��ôq�p6}|@��+�r!i5��DbF%f�'6ذ���JVȄ�=;�Nɟ����;=D��A����TD��LR�fi?�|D)d���q&��4Tp�;1~xmV��a�Goo$φ�Ӊ�щX#���;|_�b�^�bp֝�o2K�|��ғ*sډ5,��8���J�;�V�m��j�R�w��
k4����h���q�gC����[?�s�X�^�J��ɜI[A`K�B���r�=��訜g���:���N¬p���[���oWd]M#�etڞC�&;s?*�;�ϴ��.uV=YY��!q��a�(��Kl�u����*u��pUoY(� ���b�z������,�_��<&��z:���(Ĕ2m�Q3{��gT�|-h^�HF�ka�����9	/�N��W�*~πEG����O�;h�����D�]��&�<ҡD�D�%a�����k�o���{��>0A��x��R���Mv$�Z����a,�*�nG���V1s�ST�{ $\�^�Z�5��1�2m�wkO����1�-iY�Z8�E魳�[�v��'�C*ݳ�rR���T��@�ƌ���7S�ᅏx7��o>g�2�.�O��s�gy5�ݰ�aگ��E���P6��'v�M�j�Q6��ﱺ���s�	�	� �/�]�l�,-�~�_�Z/p�?���m���+�0J7<mٜn>����.Bx�'7�Y�����)M�۪���-7��ƴ��~�D�y�����uy?���P*�hщ��Ƹ8A��1��݁C�Q���'������Z������;VV�fD�,��~�xR��̢����r�����=pk�zh�"U���v���n𪎒���3m�����(���֫B����䮊����-�F��*/��t������*�!�J��}�y����r�񆅿�&(��K�mBq����ӣu��crȿa�견?sq�Ϩ3�r$�3�����.;�v���'���r���vO��+�>�`�@�5��f_����l6���ϱF����٧h�'}�n7@9��Or	�u>X���Q	&i�˘�}VJ�5� ���8�p�I�!��6+㬜�[�~P���;Y� `��6��͞��fGlI,:6߾��كz^�jq'�&���Cb8�=P��5�W��'9���z�L:��Jbп|f�$520ƛ15ũɂ_��L4��{"���aف)���u��5֯	x��L�O�A�l]B�W�����R�-�pBhmC_:��ڕy�����+(jz�J���ϫ�0��=z���x'����P<�������o���}z��@\��qN�pV�/�C�xlT�F�PFw�KX���]���v@E���9L#D2Y[�9��Kՙ�v˲��̋)+]d�����"�����ְ2��q|�Dn�hu��!��~2Um���ib˭�;_����@g�W��P�8��4n������аh������ �BpY#qN� +�]�_��F��4�፶����WoW�M�m�L�:�,��[��^��|��8��UI�lb�����K�6W��~t�K�MK���D(���&�M'�w�-����ݣQ+GZ	�vQ�AS��֘cI�'q�hO�	� &�V�/�V��K۫�(\#���e�n�!!:B<,4�n�8�%0�B n�T�����6�m��a�A�|kᤃiϜ�^� \dAZ3���cF�7�_C'c�i`������H�G
�#Ǝ�����h����b�a�[�����W���^��|��C�s)��I\��������4A��������w�jz�f
\�JPcG�.am��i�W�kӽ��'8A�U��#pg�  kAL��{�:Mj��
%�I�X:�bg���fz����G��X.��I�D]Ρ�w��5!��[�@2Z�\F%O�;�)��<�h���c?,e~�O���P���L��t��r<wSi)�6Za�]�Չq򑼍�6w��o{3�����ovG5��~X�h�p�W^	����ܼ��w���������N
�[���z��e�n8��_�0�bɇ��9��O}�]Mgq[����).�B��݅&&e�_NX�YS��՛�O_��Lw�Ѓ9s��ф�cA�]X�.����0��_f�j~��@���0�^U�
�Ә�Pkp[�֑����>ב'����9���ȈJ߾��ٴ�m);O�6/���qd(���IpJ{�)��36�k�ꏪ^���.Z�H��K�v�n�[={����� ek��V;&¥j�!G����t���n�2��j:��)?x`�T�rs�VT8!b	,q�B�4Z�\�rE
w�X���3�0If"x�"�``���;�JiD4�kD�wb�qm���|�'8��4��6w*=���	���t T�T���F�,*��j!�R�l��mM�n����(��=�L����T�V��������Y�ؠy�����;�;[1L~�^]�1ʾ��/���2�{��V9!$�E뇲{\����m�o-��%<q���0t��&x��N�6&kMw�p�g�HҌ�tt���lKC�Ũ��0R�fI�.�(j�-�9����`��A�DRK�͞/�[[t�m k�tr�>(�	�����|!��"P�x�`SPnB8qv����6�&K��R=ڭ[ϒ|d�y�铁������(┟='^�D��drq:���+���!�O��vۦJЖD��Ԍ�O1ewi6�����r��j���8�N�P�z!�!|έ=�>��5��PO:nد��p�DD+}O,��6�_��>>z�ݙ%��[I�Z��yP]j!2�N�5�L�՚�]Mɉ����nS�W2�֘>a4�q���%���o!�t�u�����^t�rt�2S�J��x����q� �Dj�Z��y.�fx�C��J�{W5Z:
f�Ν@i��0�ã�;�3��>�x|<?r{��"�=f,��g�X��%R��SU����މ�Y��j��1'��y�	�Y3nΩv~d�ql ���E{��5�7;s�Kz|�q��-��	��g]7���x����6m���,_�5Oo�e%���j��Q�x�XX�5��n˒�xaX�I5S�9ҍ���Jy�a���I���fҭ�H�(F�:'I$k9�:$�Gj�2ڢs�̜� .4�8|Df�3���Hn�Kn]sƾ�������&���͜���͐u>ױ��Nǋ�ʹ��pT]���+PN�B�0I;�.�E����5wcx<�P�b�'��,W��E۶,T��>EOp�^gVd�H�"�@{��:�RuKY2�@K�MIl��<ݞ�2�� ���c$�0��cQ`�����=��:}�a�:�����<��n�E��H�q�G�;r5����Chn]"� �O�m�Ъ�~�_1ȃ1\7�:Wx�CF���z�F3�f�k���g]';�'�$IưO��_5����������J���f#C-�A��4?�$��j��Q�b��/���v���Sy��9-br�9\ d�1f<l�]���*#�����|��x\EY���AU���<ʀua��C?�.�"�ATT�GϫQ�F!��叼�F�%�Qjh�aEhμ|���r��[=}�Ĕ��nͶ�Wa���Uؗ�H�f��r�
���~��SB�,����
;b���ܓ$(4=�?�V)$g(Z����u�ڡ�K]^po|�ڕ+���^�!��q��ei�mQK�N���Nr����йD�b���^�~jүw��W�͜�`8��O��t����/M�˷а�xՍ1K5b��=��6�NܧM=�eΊ}�_&�`h������5�0JM�Ϸ�2:ղ��y·���`���$�g�{� ���
$P�n�H�Rn�| FQ`+��J��Oe|s�T��mpbԦx����D�.~c�(��Y�Q��`�\R��e��x+[ ���G��Nx��$���P߻�� ?��{vb�UMP@e�ۄ8��k#�)�&m#p��Ͱ����6�.�+19�i
|����An�JAO���3=��ժ�^�6�"+R�&p�£��P��0+�q�D	z%F�d~A��Ӹ��m`�᠀�R����K%�� ��i�*Ny�X�G~�(x�.�d�E��%UhL�k6&\s�슲Aԯ�!+����
m��	_d�L��.VME��޲�3C�fgZ���i�<6�&Lw�Y�~1��gp�Ў�u���ќ�7�v
z$&�km�`�V�ɪy�9�\��n�]e�b�(j�0x=F�.h@ԲG�4\z�����y������/�`KY4Y�q�D�D�7uz;��i�h�^���p�u0�>+�t-�w�
J�9�K3�uFQd��.c�LK��e���%n�ٚ�����8�Xd"x��UI\sP�e|��bFq��p�ð��]�k �J���N%�;T��ء�c��/�L���0@}��!ԍʜ��V���,D�]uG3�usT�R�m��D]b�>ˊaS�b;�"a�N�b)�GP�C�Rz���� �Ox\h�G	��5m`@�L�Zz����<�f͵%�
$�cͷgɾ��A�0�hj1��A<�K�;�=�̚w{u�&���򣀧�6u�Xǈ�!�i��E��|'�>��|5M<</շ�U��;Ǖ�o��m�ìjd7�TP�H��iH6�y#�O�?���Л��:@�����Uu!O�O�+||��M�$\F�J^�}���_fOS��JA��?�CB�y��@.R���bu'�]��}�a���;�|%���"�VW�NP�;�wO�r�O�b>���#�}��
�/�^*�Z���:���6��8vy��/(��l�Q����w�]{������L����}BB�p�;�ߔ����/H:�)ޑOS��b,�|�� �{LL>x
�תMa.���gSS-]��p��2�����Y�P`� |��yGNoL7R�9���ЍG�;c�t\�H�bd����^����|�jà�o�2Έl}Kog������ֻ�sθ4�H����<�+� �nCՎ7���)�8(�&�%~k�a�3��I���npt'g
m��yeS��3}���ӊ<���x�B:�B?}^��N(��S�;�ޠ�����*[��G[B�������0j�E��>iZs�>�Qm�R�]4�ƾ�Y���^�Ϟ�}��V�zsKb�4U��_�J���RWK�1�G�Ż�Ԟc�OL(��ɪL}P�D$�{b��(Yc�^e�p��L�A��9R�� r�_\�O��8�(pLm|RQ����Ȼ�o�����|ͫY�4�+2*�iqP����ϸ�����Q�
��t�5���.�
��q������GX�Oõ�{�X�~���-�#�o�[b{֑i5����n���SsQ��0K��X��'�k��1�n��'T:��r�dh��7�w����`�7g������%j�P��y�&�.��*)�{�2�- 0�	㥚�ә���5 �q�/c�ʋ0����w�-B�m�"ֿ[ ���X��`M5�9� c�S�L�Q�����fP�+��*�B�,�|�O�A#@RA�r�in#��i�*9M��B�&�I1U���
0��m��k/u�"�u`
eR�+�8����aWZ���vK��ef��$/�ܾ4��e ���������bnPn`���}�_������{m�����b������7�s���,`��V]��?��P{qͼ2qZ���{�!\���ח��E;ټ<�q��s���M\()�4C����bx����
�K�1��z�*�s�7Y���ũ5�6	����6���|.+%�(5BO�>�UNY�<|M�s=��Nا�kpKu��,�3$���B4��Y�>��c[u7&\�V���^W&�^<������S��w�@��N�X^�t3O���DOPt�s��$�,���H��J屗!i�9Y���(Q���f����bz_��]�b��Z�tf[�K�7W�Չ}sn>��Q-]��6��$6ڠbL�m�ܔ"�TFn7���}����h`ü���a ��kX�OYVH�s�%��.	;����zś��#�������bM�\jCf� |��1�=�nyϦH�!�C遉��&���o�2m������b�1J"q8��Ac�E�P:�������v,Ӛ�2H���d*k%8~,%���\�鼍�]�c���#�z@���?��ɛ�G�����p���#:f~[s��x�K�m^:2mv�X:�G%X��!J^��z��ŭH�m9���˯���M�&	#m=�����6U���^Jx��jݼV<�q�RU���rў#���/9�蟭o��i��t*�p
��#%ct��{hIU�m-lD.!��l&����/��+�'<Ÿ��F(y$Φ��d��K���nV���F��YMU_�k�ϱ:�N%K�'Y-���=��$�Z�C���[�ӳR�~C ]>���1D��~�I{�m�+�!3�Qm�,�%!v�w����۷ƞV�.)���r�n�c�}�n�����<z�:M��ރ�5z�h�{�pi<u����ҷ"�y�L(aX�2�'Q[\����!R� ��'a)�a R��b�*K#I54�&��"�eu�}��@�o��Ⱥ��6&��n� �)|�]rPnn��r_aA#�U�&E��GC-��g��w�m�%Ӫ���@܍W�ؼ��&cx�� z��u�J����!�88���G�L=�h�*=`�2O�� w윻��k��/��I~;
��O��>�E���N��U�`���Ə6m"���NW1��t\yx�,P�s��INǾ��#�'�Nv�SM���T���^�&4�K�Zو����C��2�*
e���-�S
���Qz��$�!�������o��bv�]Cg�9�m��TI�3I���̝�F� �j�@u
�sY��d�:�������D�/��D�z�,�� QW\Ft��9�@��&�nb�헪[K��W�m��(_�Z<[��;�\m��Ha�ߒSzӳ.��_2�\'�����_���l\Ak�ouu��m�4����?X����@���&�&���ն�Kk�4�i�qG��3����c�UB��t�-�Қ����!A��UI���pyy�8p�`���d��(���Jяg�6i�d4'��G��vR�Ө����J5H��b�UV���˃��@��6�b3G"YY7�3T[�,?i�\�%b����7)$	U��w76�_7��ɺn���l@�D����FZJ O�݌М�hs�˸�qG��;�� ���}�#v&
���5 ����5!^�շ�C;�	�s����1m�a\����	���bކ�����y5�3�!HW�1;[�,�j�8�O}�b���=I��g駯Cҍ��U]n�( y�7s���_q�/=ԧ���jMl�k��Ҝ0��N�j�+JK���Zc�HO��,WW�1	�`��G�����q=�1�_��G/T9-�-��ӥs�,�*��4��B4YJoG�R۶[x�S!�ج�R �N��T;�D�ӲCdR!��-���9�Q�lm?
0�,5*�M�y�9�����L�K�<��T��ra��)"|��Φ�`����R��f��I޿��ԄQ���%��e�+3�����5I�i��"��r�q��W=V3"j�F�r�j�*�X�'ܬ6	\lg�i�L��:<�Og��2s�H̝;k�)��ɺ��RQp{ʌMAü;d�t�>�(T �^@Y���!��vm�� <-�������PF�ܽlq�է�0d�hN�op���@\�f=�5ۙ�����T]�Q�Pv����n����mp�r5Ug�$��Z���<����'�&t4����N��r�$x}�Z;���&&0Li;�b+ˤg���k��y_�i�&����V�Q���Y��A��P��N��G�K	�C��LL�8u�N`h�=�#`,0[K�*���^�'��(�~$��$���`k_��g_oU;�� Bd�-��,l��&x+Rw�V(p��Nϣ��V�d�M[�i��"��ʮ=�p)���~�F�NC���'m��f�;"�D;3�Ii�����8�L|�q@' Ծ'��������(i�5-�@޸haT_�"���]��9��+hS�UN#����j�ʿ��$��F��v��o����(����t�U'�����+�Q�#ۊ������x�/��N)V/f������ӭ��t�OZ��e+�ب������?x�B5���7t�&i��7���g�1\�(�9�̼��-��R�d=Х�!��(W/V�UG��x"�Mј��I0�V���։�	�-.ȖߒX��jX�HG"�ju�y�� ��>i�t�ʒ�H���Ӎ�e�)���N�<H_���G��s����Q��n]4ϟ>�8:��:�����L�<�'n\��R�}+���1�?�R�R���rU0��N-�1;�����] ػʹf��I��#�C�_-��_�j�sشd���w�"�i>�3��yp�.#-�%�ȵ� ���N�5�M����~6}彙�o�C*��,@������M`��^2-c������v$�$�d�\kz���eFV�]'5m;�z?�y$�V/#�q�͈��	��ܲ��@�M_z���$h� #�.w�5��/���6��q�-60@V�hP���y*�Mڵ��X�X�p�HV�6��#/pFY����`S^�G��[�!�2�S� K��j���� [�<���%HW�+Yِ!g2<6�E���m����5�%���������4����f��t�^r����������	c�6����6j�$
d�O����=�P�p�� � ����ւ(d�qwt}.:=Į�Az1;*&yƚ�'�]�����-�b.��稼�S�F=���w���{�ck�x���l�C�8翍�%h���:���4Si$�c|�1�>�b�]�����u�Y�Z�B{�{"�N�(�
��uV,�P,&�4�~��QE-X*-��4.��/?
�JA%=>Hw�9ő�`Q���t-X^���:ݠ��z5yOr��Z�k��W�X��6�L��r�\�w�y�����!B�	~x�_�J|�b
�����s��m�x����*5�LS���15D��O�4��Q#��а�_e���}e�����bl�J�g >v`�>���0�ǯ+�{� ǜu������aC/�{���ވ�?�b��@�k��]������o�j_��`pP�p��P@-��T�5�\���y���a��L����x\(��[�,_{D��݋� �'� U�)>�"�6�4��w�Hl�����@�p��`dtx�!_��������>���K[;(#�A�HJ��-	�b ظI�����K���J7�v
����<!G<{�|���{�,i2���kzB�TuW:�ƭ��L��Z@����E�.Y�آ�B��
��:@�ճh����Y��ޫ'�{�5�{�*�λ�Q$`ذ�U�1����"�$�ic�Sj��jѺ{=_mT@u\�t)bU��h���v�I�6nةm�E�Ox����U[Z�]����|�����I�-^ȹξ7�1_}����R�B�6Z�g�_LT�$��Y�,�*� ~��xP���z�)�.C��lB�Q��8}f�z�2���C[��o���^#σF��y��5%l63�]�CHL_��v�K�e�s����&!f)�J�י�}j�P!@_��(Bf�CHz���	1��-��A���m��!1w����p�3���U_�T��g�0��'�O�m}���*�sz2/����i�Ǐ<oͧ-�ڛr��6���1
�����
�U����~�0�h��P���Y%"T���S��Fb����v��_�B�]5�Ը.7Ph�����T�7��<�y�%�wR[��J�Q�.*@7r���Y�pN`�#4�J�}w`a> �m� �S�Ύ�A:Ѣ��]��f.�#R+�V��o�p��sSm�3�R*�H[��'������������w���)����?+W�{�O���Z��O�"��`8pj%�@ݩ5]+��w����a�"w�9`́d���Á�H���q�zM�v�l��Qzq6��V�����O��H8����\Y�&n��J�����e���y��!C^X���_��$��y�1A+G��,=J� b�>`���|��=��yΏ�L'O���O�ȶ�!�h0SL��E�B�%m�=�����
�X���7��|F��xW���i�n����b��������Գ
-�����`[ϛQ�7�ft�7#H}�v��b$�V>����e�+�DS�O���=]�NW�?�L�l����G1K�,�>���G��B�G<t�m5��P[��$��+f���v�ᬨ�t��O��N�m�3h� btA���1���r^��I�.JI4P(�"S�^�|>�9�hn|
3"�7��C;�*#�	'%�C%�n�1�!.i��o��g���{4.y�,�|,yr$��?V3BA�C�}s�M���y��ؠ�}vĩ:^���n<�w��u*	�J�z�������������ԩ~���H-��x׽'m�!Ī�7���Ko˪Yo(�\��q��+ǜ���X|X?���DS����@���a�~���^�&J��t!�����9ѹ��������#ʵ"�k"Ц�K�"��}�}���� �GN+�R-�zmM-��P-��X�_���;�C�*<�\Q'&�}^��z����_�4��ԇ1^�t��f�!�U���������g�d+t��=J�چ��J��b�6�Q���1/����(�k��2BV�V��䶙�z��S��"F�K�g���2&�=X�d(����̈�w'u�|L�R#F�Ի�^_�u�@���
�f�>u�mr%	���,�����ĩ��S�] ZJ`RQ|�B��'7�������'�(4
W�Go���1Y^@�o6wt+v��:J��=���;GZ��>[�����9g��nGڸF [`1��1���I��iKn�S�M#���f4��z��|�R��f'��A�IA-���p�(�{�@V
�\E�G!��vfK�v����lڒEύ23H�$*�q�����M��*PvG���s/۰��+�=u��:%�L��-�#��}3x`gʊ��.Cm��� B���"��H܂�7�%���hH@�����/��1�5�ת�o�U	��Gu�[�JdZ��4!%Q�[ ���&����yUP�6�d���(x�(�N�L؈{���a@-�dsXh>��!��.џ<>�0ٝ�hàF�¬b��ޮ��0�<����M��W=rH5ͷ�NN�����7�l��z�&Qh{7;�6�[����d����Vx�a`�(=����o�{�Bw}g^�dt�VU	�Y6n�\���+���t����&r�Nl����ؓ+=��rau
��<����h���_|?��d�2P�]�p���j��e���II�x[47�X=��ܦ�����5���b�_-B
��g����"{Tb�:i������^��	�4��t&���1�G�,l��\��E >���s���F��.�&pk�{NH�^�q��-��cx���j!%�	"�ȋ��ɧ�c�|"�������9m��K�%�#���)���/���ċ-ͻ ���S���o9pwuv�>�_c���maWR^��@M�xF�q״��U{��)"~(��ԮZAbiȨ ����R�!���
�y"f�;�m^����k��o�C�*�ʙ	��s󶳍)��lX�G�
]�T����YIr�{�/<b�sE�{���,$��H��]�w�������3���U)����K�hR$�@�&�-�X��0<�������� ����@k�� ���<xy�w$�i����^�gȩ��;�C�3���޷J����/i�$̍��u�Sj�D�q��ovl���	�}�/7۾���h��{ h4�Y ��C���J�9{Z��-�`�^�Y�p�G�2��XDS�O{�rm���'�$�����m�������DSMm�J��s/��H^�e/
���.Q�K�3@�Æ~>�LZ��
2�tk �c*�/G�)���#��d_�b�X�Y���h#�F̈́���M#�:K�hkɉr2�|]W|f_�D, *f0>��I�b�j�Q���=?6�2��P���0 7�A�.�5j�!I ��^�=x���Ka�9/�C~H(JO�*#�TYx�,BrZۦI�H�]v������83,�\M�ݶ�>��F��E��6��U˜��g�8l��F��5�eC����[�"���p�B�G�A��F��dH8��O�����?ޑ
E��ԛ�?Q���\|�3�����a�yD:p�|3��T@��Pǟ��rg��4�H����ݟ���}$ù�%�BcܘF�f8Ű��-R�8j��wy�/Y�(��� ���`{��\}��n��}+X��ݲ�K~�c҅tуb��ҧ�g#��ҭ�^"Z��FU�V�Ѣo���ֿٝݽ�n�f�*�@a1��7�ܪ�)�2�ʝ32�-~`�����8�}}��0��e7�d3o(�0��]�j��I���c��$I�cAG\��|��%�I�5#�@�rK��R3vj�+�`�en�T��;�5�>ɇF?M3SY��Wk����@��FƜS�=u2M��PLO�YPG��
��d�ۋ�� ���KCU��{�UF�����Ρ-v.�k�s"���#z��hJ�^c���	����v�/��|ʅp�;wlx����R�.�C��u���&���'G�`3J���,��4}s��RG���A�&���ߚb�N
�,�s�^�J�s�?�y�EwNUյ��85r�p��z��
���$���k������fxJ�R��HW� -5ckGd9�̊�N}�b��'�����<��_�����?5�F�E*N���\�߉��6[�<�)Y�k�����F_��:�a�O�;��~�N*.A���
2}��x��4��'�vTU��jSS6���-��^�A��M�|�?� H��@�OY�1g�;�v��.��Y���3
���I[%h�F��m��	���QO/P����X_�p����)���XAn!�e�`-�Q���TD��fU(c6�
��`y�?բ���X`.� +�����/ny&�eg�a����(ҋY�Vq��hw����gJ���~]�i����UD���Id���A6�I~��qn��@�]����[���s=�x�7��W>I\�bX�D[n0�u�4�p��Y� �J43h�7Hlbq�t7.����C��"�k8X��P��A���=?������j?P=��,��|��7f�^㏜ʡ� ��BGZ	'��k�̎A-��&���Z��H�����.l�"ī�E�;���� Ճ��X��l���3�f�?�0~ �Ǡ��r�hc��%��O&��?��wY�oJ�b:���3���DX�!�2ܚ�ͻ!i�g�� ��%���S���4��ɜ?B��IK-ǳ
W�p͜�7�~d��:�(ZûsDw�Qb��6&�XvEP�CY�j��/KA�:���p�Ă��q��
� /�)¿f�(^`C��E�A2YS�-�G`;���\���[�5"_S��a�ڌ��&!�We?��D����U-m�xM�:t��G�Qz͡ʞ��`Ոv[O���_jw�|-8��y���{�oѱ���dEXڣ���&���1�a6��B��;�ٗ�Py1��]�FP�N�2�"�'��ʊ���I�kC�\ㅊ/��Y�Y�&��uK��4�J��*K����鎄d���N�P޴�=u��?Πw�_^�c���xպL��^hQ"��U�Ӧ�|�K����׷�nlsM�6*�����.��"v��X�ۆ�DC��{�C�#9�j�F타`B����*�� <����O�!�\�L��ӿ�Ֆ���;��*�Y�M���k��/>�8�]`BΎ<�x�v�[�l�,
������?}�*�P��x?����<�����z��d�i<k>��������"ڀ35���F�Y�wﰽ����T��5�l�e�2Yנ����[~��i��^�������Y�%}�W=�<����d��]
�d������M���g6�c�v��>6��}�WpI ��n-�y/�O^�]��;��[�����2Ք3�����}2Q�'uH8.��E:6nx�@�PLo܂ύ<C�<����s�u�]���~��;l�$9��k��@	Q�������jJ�T��h"g��.8S����Ƞ�o��T�ЌX5��}�������S�Iʱ�w	��c12-褺��x=>Dk3��p���kU�G9�M�̆`g�b��Z�uݢ�'��xI�I�"����LĞN��\ܪR@�lh/��4w�w�ZJƟ�
����3l�-&���6[j�7��k5nYS��kf��	�s������
Z���x�K�2g����9�:o�*� >�Q��Gp#�|�{��u�q$��],�� &���D�:X�?H�_��ߗ�H蓷���P�'�g�y���l巟ѽ��'�j��Ӧ7�'��~S�y�·D������(M��	� �ߤ��^#ɻ��&kX�2��F�	yr�l�f�����5�#���(ym�yPK�`Uk����o�d�!`$�/�k���y���b�v�IM�LX��f�K�I�Uz]Fr��#@Q`�!�xY��N����ĐZ[�����!Wfn�׀4:�H�+��3��{��9�X;��|����ڄ݀�'#��s:��<�ݐh�n�zHj�/YY����s��\�?$�Q�Y�_���5�gUN���Yr�w���+|�	[/H
���� 8��l���~�*�i����ɍfn�~tj���cQ@w#j�{�3�S<�t�)=3v��Ӳ�m��+8�Bפ�I��uٛ4Qv#lj�{4&%=�X��1�X�u�0���ڋa�C��,����Tu��p�җ;Q��_�Z���8^iv��SC@�
��
*��'��$��z9�|��y���-��d�.�d��^�ud� zSbg��ɧ흜<�����\��+_SE!O��	�=[�
>�jc��3�2�*��r��]@���v����5�����*Q\������)��,&��얓����	�>b"�?� 3�����Bk���Λ�m%��^����L���X�Du�AA��7l/�Ϯ)����ֈ>z��ǭ,�XXr�;���m#Q���(:�r�E���Q#�$:����rn!��6����w�籧���S��yMq/�$�K������[T�>�G��d�����ќ����W�ޖ�1�Ap�N���C�D�`�������;�)��l�X�ˆ�#�{h"+?����쎝���'�R�V��}�@L{!��҆�v)wϩ9�g4�dI;�漯��^�O�:~�P��=5g~�� �����H���
��Y�W�W�4�:�����q�mHǛ���V��>`f�'̐��_��v�tQ�~S�nf*�1,R�ʕ<�3z�fӯÊ�>fP(e�$g���e��#���
�d�,�͔�O��lܘ�(��x��W7��H�������~��1F�(H���*.���`fR !p͂��i"^m�_b��j'#!�2�
G^?rys�Jy�s���2B�S3ލ�6!����l?��׻&`~)�K@��+ V�j��2(3��ڑ�@���,f��r��0)c����7hhe��]�����]R\%.��r&��)�Y��Ry5�\k@S ���ޜ�����6u��H<g�$䐮ib&�Zd/ιPi��9Ι,յ|+˯�ЈW�bt����#���(|����g�H�P^�4��P
F�9 ����w��D[?&���E�8W.%���a�с�Z�z:�u�a�6��wa$L(�ξ��1��=�[_b�.BLu?3��$�,6i��m��tyU�!�K7�"��W潖��)M
ZBc F`@{�٘��6�z÷&����l>��qN��?Y".]`x�f�6�7�7C 폋ʟG\Y���a6,<��%о�a�鮀xk/]��>�O�76yYy�Rm9i ��B޼OԀ΁��������2K
��Ζ��-e�����]�f���|0?�ϱ������{�[]��7��*�/[QN5L�)p[���r�����P�ေ��R�'t��&L��#~A�rŚ�rb%r���Ft�=���>��L���v�7ա�Z8��M�/H��L�	��g#�,�I���������UW:{Q�ȨL������r�ժ{�:թo� �A#m+��AO��� {`�C�5�͗,:̀4��{��Y�n	cJ��pR|Oz�����ߑتec�=�oj���-�E`)|�'{~i����O�Ԑ�p�Y��)�ٌX�^�mD,}�a���c��䞆�UB�|5�����d�(T���ݷw�M
�Yjă�7��s��-7�b����Bw��F�P{;����0u��ҡ�f�`١j��yv�~�L]�q�wѵȗ��bVڕX���	���V��C�X�0d��*m+(�H�RC�F!{Vw~���e�{�l��̣y�-:��	H]sm@��J$Hr�U;�W�W\����GV�sl�ށ��<���2%����3+��sO�6y*<� �}�n�J_�f���|P����~L�u垏�a$e&��8q��r�b$�ю�T�$}J����H�P�h��b,���^A賉�\���<ȷ2������Xz��-U���Vk�ơp2w����L���ۤC�T5�Mϟ����#�L��%���4`�E߳RO�l��s y��d��QUݹ^&�u�*c�U2T�{��ۘ(N��������o�t�d���{�QњFP�����=�Kn�z�,��yeJ��E�T{�n.�	��j*��洡㟮D������<E�Ͱ�H��,Q��jh"�@����P�������XR�t�=W�^w�UT�Ʌ[�u\��mJ�/���'�G���ď������7Ϙ�N�'1g0����0VP�h�Z��vA{��諑���"��m��q��0��]� �8�!P�BV�*#{ºLF{�L�#��}��f��q�:��B����6����F|���Ve-}�&񠜛��a�3�!��o��!����r8)��B��-V\�������ߖ����7��,0 +[�Ǔ)�%�%|Z��<
n5�%��p�1ЅotI�_
�������I:����ҊO���P&��K���		w���B1� �w�����%�����Đ�JZa���$`fO6�������[4@K� ��/��Ab5Y��zZ��7v���G�̬�z��#�_�����C�9�&�V�+p����{Ѩ̀�1X��f��,O����������.�;Za�7c@�(�щg��;>Q�<�}��ljf��tt�<����X���+Z�m���H�G�mt��<8�~���(H9��BToxX,R0زp��OM>g�*��rA�Y���s�x���f&�z*�ߧ:�{�GC�^]���e.�x\{�k+0�ކ�����聏���;������'Ǌ�������3�j��;/)ܞIXz��a$m=�;j����ʳFN{9��,,�/�BhP9������ ��L?qPɱY�����=ןH�Qb�����Qj�)�H�vk�Q8E�����Ј�o���z/G*n`pJ����x���_&��B!��?����uh�x4����-�cC?���k��V��f�Ʈv������bi�iC�,�'��B*�j�Oq]����u�P��H�l�7��ޅ��yۦ}�J�!��b0�׫*���Lr�w�)>Qg����p����󬔕��O\-an|��	w�(Ԭ
�z�>! a ���U 1ލ���n��t�7Q
Iw=���{
��]��Z��S�ɩ�A��X՜��r�<��t�-.z5U�G1A2l%����7���J�\0��^`����H�� ΅I���<�OG �?r	��h�I5ϛWȶ�僜B Bz�b:�#��� >�6Yog����n��^>�G�c������p��m�F����iwZt��2g�z%=�I]m�,�Q�Y����Mfߓ��WI������g$vm��LL�U��]��#=���ζ� 0g]�2U�61���y��wf�:��k'�T9@&�����D����+��G\��Of0`"PN"�)ӵ�D�)�l��5v	��yI�1eP7BE
�0ɶW.���I�"��H]>����ٛ[��r_�R�z���$�X�˚:ٗ�_�X��s�F��Xi��R���c��	�<�b_�]�Yw1�[�r��^{����D:�u3#M�>.��М��;�N�:]�a�M���z���܅���	�T��๶���i�dsh��2vm&��F�o�f5�G| F<��-���zZ$�4Z���d��"
a���_~P�ݖҟ������5�J�#{��𹕊�Ȯ!�QV�J�.�+� ���Iʀ7�.��ҹ�d��󦔁3E�4Ǜh��[����4����nb�q��3S���EKݟۦ�82#z�U�2�/m���hJ�O�V���[�_穐�Srad��&*1�vq�?"	�I�L�$d�5
���Q��Oa��L���G�$�h$�)h�V�|�ʜ�'�E��o�@�Z�B#$�R7�S���(TXW��6�69[A,`*���àK�"�j9�8�o��NcW?>nb�J�W�=icl�\5��� J�~�٫��M�х�5�C<?��;��1�{�͡"��X��l��:�P�+Cs�*,X�.|t����o���c�K���~��W����ԥ�s`LVso[eB��U+�%n�f/?pn~��=� ��v�Ѝ�����XWX�G4����)#�T�Z��FZW?Yv'�t{��%.��-<=j��y�����s�ڞv�p@ʩc� UX�!�r�̏$?�Ǩ�VK��5��x�{R�֠K�	m�؞S�d��;b�'|N����"	�۱�ͭ�S���(@C�f�h*�g�dL� �"(�L�PW���I�$�<R�RԾ�&�$d<��냪g`�刯��GW�%L@
�y��ų"����lI����+p�WSF_,�� r����Q�vno� (J�F�S>@�*��E�Ƅ��v������`��7��w�<V�"�b��O��!L��p��?�iX�)!@�g�a��Z}IbnL�£F˧���~Af2���/��u =��� B>)|�%�OWITo�˱�EF�}�g���>��9�-:T�u�W��7H�H:F�������J�T�R� ��Vu-c��Z	Ɨp�UK�e��x��������vuNs7�ՠ��ȥt��&�-n��#cCy. J����~��IϤ�i�
@�M���#�'Qb�䑜q"��&���%� #�M���8� ���p�7�HX,�d���+��H�ب|f��vYp$QT-pBE��q.��"ĩa��Vi��I�W�վ)J�YjX!-`�)�ǵ�C��i��1C#�d
�t�,�!�qn¯d�q�-�;}N�mE�`4��=����xZM�.��������{9�[<�G1�+��,M���^��ӹ��=zI����I真 ��c\G�s�G�^W�@�0���s��_&4.�j���du�`4N��/�ÿ�����v89?Dk�<�b%�#؏���$}��.is�I��O+��g9kF=^U��}��/*h������B�C���2̡c�=�E��|���Uǌ�|�5��u����1� \�k���Dj�T�v_�����+��B=����ski2ǰ^��9�xfBՙyH_#p��k�
]��/�'_�-�է�Xq����ŧlM��I��;��5�B����D|g��^�k�l�9��ՆV��L�ej���v����|!w��E k�5B/�BC�*�$��4�%xKo/�>��L��ʾ�V2���xǤU��"��V��fޑ�o�!�M�;O5$��l��֑1�ɍH�_�.+I�J}H֍��kE(tn 	������vB��Ү��x&̀1g��u:�1�v]��܁;y����u;^��ӽ�>�ߋ���� '犯��h5.`J��0�:�����ykF�iv4���!��½D:�D�V����@�l�3k�6-���ޞH�C#��:2C�ʀM\r
�8Gq*�9����V��z���Vp!��[��)������
�k�H�1�x(^��̥J9o,H�^��:8+kGl�%�4�\qI�ǳj���:U��G&��v��>5����e�e�*%E���Y(-�_�G,�\<_�-�]���(�FÔ
e�\~��#Ζ��͡��=7���N���k�����0���Я�t�i�1ʔL����]��<��l�m����!�#��D�:�y)��䓄����v���a�3�i�<����6�^��C7�D��!F�M1^��w<�c|�	�`p��7��s0�(�w�B����Y��+����{�T�T{��/:o��޹9�p��S���0�
�9@�Eq�x&����b?��{�q���5ּ�R�rH���5	�%����R���`����s��3�q=j��]����ʺ��o���w����;,���6-�;o=��2�����~-���'�C~! ^�B��fI����hT� !��j����&,�)�3�obj?
�WA�5|���ͺ��s�X��� �e�V3?�r�y�u�i+��>-�4��_���=��=��aa��x�fQ+`>qk�X#`��q1ݹF�z��g���t �����Z���e=h��G�甀OI�g#?���6�N���A��d�\�`��5�'�|�D�b݄�����'�4�#1O��m=���1�S �-;T�����K2�}�ώTWo�ΉR+�����.�aQv�5@0�?���a��H�]Ю���a�����)D��m����3��#֭����� �����7ȕ"�.� K�P6~'r�U`d���@6%�a��b�/�<i��jL��	���=#(�C�U�k*�>).j�2�ҴJ��
QRG9��䴡�?-��a��>^gq�K�������+�(��B����#�2Z�{�b�*�����s�4i�_9��Ԥ��e���0Z��Q����)��O Zu@��/n�����Ƣ�y����Q�'l�*!fT��(��p�7P;����cC�g!x��vڀ��	�6B)��|���G��D��Q��ķ�0/�#?����Ey�o�tޝ��u��\&s�4µk��߱�]278�n&�h�u$���d5�1M!vk	i�u�p���k��������3�.�F�;9A�[��Z�+<���@$�����]'���x 0��;�)kGD��r�۟��4E��~s9�ŉC���m��<*�!&�f�g�?�)�E6�2��7H�Ǯ�E$�8}�C��@��[�L���vNgZ��v5��S5�;�
��`3���9m��_�ɦC�X�p�� ��+[�T��{5-'��͔�5W��`:Oyb:|���ȩyA�x����oݥ3r`��0�w"�o$��V?ĲV�����Տ�������:�R����ӱ�(�|~�z��P���(=7*�l5����g�c}�B��f��r��;)�+�h�tW��}�zzn�\�\?D;l���2ir�VkLwx�5����|T�xb��D-�Z���m�=m9{p]�݌vMkՏ���2\�v��?�1��D���ۇ����Q���؂=�M�%��+.D��n"U-rs�ĲJږ�t���*6_c�H��IW�8<��~U<������"��O�E_��p&�scD��	s��S'_ȹq�AC�L���z1�H��?����m�� O�"����Vl46��u�1a]��I�[3� �xϭi����7�������nw�ǶI�ƍt|����ӸQ�����`>�0����Y<��"��;�� ^�u�/�B 1���$;�)L�'�^|��_.c.�,c�}��.�Ǯv^��bHqX��'j0�q� ;u�h`�0��#���-\�wq���.�Dz\=�����l��F�D��-��+��+����]�Q�ZVC� %��J��������7�����J��%Ɣ�y��vĕN�f��叄	v�������%�R@v	���@{0,�3��k�*�s_����:�:�6��aE���v�(���"*�<��CD�1�;IP�X�E�%7����m����z�;Jy�
���������S��5�J��H1t�2��Ȃ��ܨ�5�?�w����,1	�����Qj��˃�$�Z�:_%�#�41[{b���1�����B:N�v-�Fȏ�}+�l���-ӔV����3��.��}>1/�Ä�3tez<�Ĩ[�x=v�Ʀ#���&��ھ�l��*�^q0~.H��&M�����;��OSI��Ω�&��V�d �6���|���Y����Cdt�����w��7�r�=�c�G��:"W)<

"�g/��R_3rM6�ȽQ���e��E��X��pԚ�1�{y����P�E�J�WWZpV�d�ekN\��P��ƴ0��È����C�e��������N�����)bJ3|�R�W�y:s��WF����&�"�H�p��{G- ��P�,�LE����k��J��u��A�@�RM2e�Cs���B_նy��;��
ܔ,�e�}׵�4U�{�y��mq{�{�,Y��.�:��j�c��'*� 4ø�˟�Ǥ# .�Q�S�V��(���9��/���`�p�V�PS#m�qG�����J�_�1p(��E⊨%�M��!D�* ��.��johu̲���d0Ωw:�d[�h�[�-���a����ځ��G�ڿݩ�I���GqV��\45E��{Y��HP�;h�r�^م�Q�+kLGq5R�g�����?���9�_��W�VUĴ����I~>��������;����xؑE����T��C��3[b�bm�IJՏNV�XB��XU��Fȩ��BI(T^̈a>���;
̿Ea�*��V�wy������
���Z��[�VZ����l^2%-^6�ԧ��)#�FM��wZi��R��^wLʗ���w�Sl�⫻��l!�V����8%������S5@�vA��:�R�!WjcyI��uL��I��#�s	�1iW�{��;Z
5�#��3�n�w$�2�&���I�Ѥ)r;�i�3=X+m��ܮ�C����*����1��LBHYl�����瞠�"Y��$��_>D����{�v��akZI�vm�p��)�0��g�b��璣���f�s��B� �4g ����4�W��0�HG=�c,�|�X�F`� 4ȣTӌyc����3L`23V�/kG�-;���4�/�e���-OX���#�]����I��/��"������e�͜s>Y5�~y�SJhlI������@�mY�P�r�FK�6����˴�X��EE������4Y��W�`�#������rD�w,�o�$�w�x�H�s+iQB���C���2;$��CE+}��%p�1��/oD�tVَ����O#6C�e󙆼�q���6����VA|{F(�g�u��� )�B'C⡊��c����>Z�3�o#3w�I��'~e���˂�Fd��>�j^��I	x��<��Vy�Obt���P`XIh/1����s��t�Dg��򃮎l���Y��h0 	�[JҐ��@�\w����D�����=���������v���6�/�ҥ��3C�G��UI�������,�:��?~�Ù�֍�;q�f�)
L/ 2����z�� s�ρ}������zj=e�Q�z�D�qT�d5�sĞ����1b<�<ϜYI��I3���h�sm��?��a�
��>�f�������$Y�����ej��^ѧ�Q�������Sq�1�)]�ʚ��*[�r6�6V��f8���[P�����̸�6�j�������ಪ`��tCyҞ��E�I��G��p���Ѝթ�Ύ
�!�I��)*׷+P�w�1�*z�}��c���a��S�[r�)
J��c���H�y5�\���^�q���.���w�v�]����q�nQ���J���>���V$J����G�%9{q��A�_�j�R��f���|̬z_!���g�����9TFl�
��='�2<l��B���;xXkC�g3]I��;5tν�����_ ՞o�r_Ҋ*Ӷ���V�Qd ���P�-]2E�w߄gc�y5�fy����. |�c�H���C��o��n�i���ZL��pZ�7�b^蒍���;R�N�cb�3Ƃ9fu/	��[ҿP7�1�ѹ��m&��s���8�2���վW�w-I�V�-�}$-y��z�ȩ~����A��.W1o%�q��Q�G���X�-*^7�}��c�g]{�W7���a��T�#r�$�5��X���̞�#�-����_�s��pb@�+&_K!&%6���4f�G4���=	�S6|M[FAPp?<ь�������:��� ]�??�A�<b�jjΠ��b�"����Ͼ�5��c�i�:�<֭|vQU�}>"i�%v	���~�Y̼�2��?��h�|�9A����4�q/����s�S�6��bʳ�*�[�q���,��}ø�����!��ܬ3e��aμA�����j0��Q����^/�ǳߵud�7�������e�ǽ��7�}��S*j����.zW-��#�QCO�Ѥ6E Y��e���{�r+c��c��s3�:�H��DW k���ˣ����e���yz�9f�ؠi��0M�եi��{n��|��d{2�b���̪��5���r@�P�	���xO9�cz���3ŏ�o+>�!ןz'�\��Ӫ'�F�sxy;a�� 6���[�A�4���`�����b��~�[���6�r�\8�l=9!
?)b��VǆdW�&��&��m��;ٛ]��G���� k�^�[$9N�6��Q��aŲ>��6��y��Ŵ�#�_F�Cji:�l��U���Z��fa��������Q����伦4�1���\0���T��=���"9 �1�Z�����͢�#\��+���FQ����Ϫ�LV��Ј���s�%ؗ��p>�`	kxA�+�LɊd�I�.�V��.)��t>S_}v�	�so����ft�]�/��V���g�4�qt�!_��3��@��bh1��l'�B8�
���C}��kp5���z_�q1B�&?ǡXn%U+Ԟ�1���%Gk�L�Ŏ�R�ϳ�����L��ň�R*��ڏ��\Y�yA�>��IE���ܣ`NX��Yu��5�����;�ģ6sLp��jM==�f�e%<�1+���f��1+�dN<E>�]�&lr�n��>�����5�o�*�0�Α���YN�����wJ�8y��-�k�g��yY,�4~B�#lcU[�F�l{{�0s���<F8�,D��0�5� �Q^��|�_�2�3P����1�J�ޓ���/ܲ皀C�*�_�Zh�h�F!�^�5��蕆��Ȁ%����$�j
���wS@]���SW����;�����IU�����k�	+����[z��d[=�>g��� bK��&V�fԢ@\��O�O�� ��%�*�c
��Ixv��*
t�+<��+ͮ��' �����_n8��������+3>/�Ǎ� �^�(�N� JGwA��Q�Nע<�Q�jObUM�Mq1K.ƕ0שYr����ӆO�Fn]n�f�VO�w菨e˿�e�F��
����q/}eT���t����AJ2�Y��e��!��]p���W�>�(��-�Q}0�m�O}nf+xV����5�}1��ނ>ࢭU*�>w�9`V�{)�{�.6C]�$�l��w��N#0[��-uKYdJ�L��l�n������	�D7[I}Ni��O �]rV��ˁ���;���>Ɛn�	���P�ݨء�/����Z^TOL���g$�$���=r��n3� "���8��]f7t���C<��W�	�A~IN�ѣT�.��	�"������z�c���!Ȁ�Ů�8X�ꤨ�rXT�;魃W��A�\���ӣ$~C�y��C7�M"x8�����zM��j_���Ɍ<�IPN߽܂���T�~@���8����#�,�[j.���$��X� �w�63�t��L�3�t�I3�ukl�	Z��߽X�*�B��y��!?���?�}��i��R%8��,�����iFI{c�P.&�}bͰ!��!/.�.?��X��Y��9�q�x��8+Ħ�I��3���,Fq�f�F�&��ߕ�o1i,~<jg�i�{>ն�_��������`������s7�j}�mE�+�%ϐ���&�J"mv�������j�>��Nu�`�Y�x6ؾ-z����+�B���`3:�����6+��u�J�U��5+%*���/f�(�U�����f�������OE��{��]�č���AU�9��˗���Л;��j��2��gew��\�$M����=]� .�Ӆ�6�����u��l�m+9ܗ5k���A��z�~�e{�]�Y�8Z���G�,��=�#�:mb�5���A�#J7���M����Rc�x���w������y1��c�ˍy��t�|_:Sخ���'�ȇ���g�%��a��T���9OZ��YE v��D84�4h��Lc��u`Ѝ�&�xiD���)�1g�F�Q�������i�`n7�K�Ch��w^�1`=�=�b��7��?2�]�,�or��;��~�����#�z\�Au������\�"f^FM����ؕ�#�Cc�h5�85���OiS�稄:�nu�j�q���a�9���G�F�c����jMy��×Fz���t�;� ]&���KQA5!��p�Iݣ(6�>_�+L�C_�w"q�S�:�����/�ʨ�L�!���=��[��^&�*��3���Ci���-q�BNEC�.<p$ͭ������][E L���t��Xm�C8��v!,e��uz�$ψ�X�K�t�!�g}��*U��8�DzH�;vr�����7�gP���N�eF�똡�K�DE>7�p�.S��M���)�۸��\?��Ա�Zh�?�I�q���~Yut�q�+I_�}���v!��:NU����Ο�������:ޢ7�Eށ�<
;lrH���b!X�����J#�ʚ`��B%�۹12��3��j7$~�*�B��	I��_��Ğ>����Χװ��ԣ�Z	�g�%�m������~i)���z�Փڒأ�BC�$	����P#��ŧ3�F�ƯD�k��]�1�3p'u�y#�KH�ʀd����j��������8�P7s8�б](ox��]�(Wb|�3^)$$n���+�$�nҲ�h��e&�@�kl[��F���� ����o<y@�gR������Z��p�8�C�T.�z��~$,��<��n.�� \ ���4���*<~�]Z���φ���S4�L�ȿ� �s��Ix���NͷT��愠RU��%h����1���P�5����B7y���%h���ģ���
��l��]� ��,O8��8PN���``��h�I�+�ک������I>W/Ȏ>�7��,t.s1��|�Dwk�(#���FNT��B�e��}liu#�[O䩳F��j6����t����!h�-�s��F�%�WE�j{Z-���ߎud݉keҤ(��C��}Kz��sT!%?�r��w:zo����3��@�*HU���0<{��j�����e���f�:7�q��7�k�v��
�����F]��Ib�78��1j ��nc�#;�9Oo��P!h������ [-��W'{��^��BR��8�Y �s'�&tz�Fz��Mف sJaXH�i۱�A�Hp�>;Z�V�N���ʫ�dq�Oҥ@�B ��Z�;v���ƪf匄�S�����W���˄�h��sHي�I����\�"���&��^8-����Zq�7�n��\#�L����SrE7A�0�$")�]�3���)f��Cp)�:�c���tI�ZFB�j�@��E&��� V��/H5Rq���\�������ޗ6&�4�:ˏY�%4/'L�T W}��!���'v�i���ȧ�E���*��D����|��q�y�m��G��W��&�|/�&�{7�A����=����%D��p�KѶ�K<�ۄ4��t*��>5��}�R�����/�_��jAK�r�@�R,r�n�}��>s紿�*/>��`��X�!<Y:<�1ԩ!r����O���=�Q,�4��q�������<��"s��ѐ��4c]��G�O�x�Bvz*���A9�a��]��ʔ��R���#��>,��<�3���%F �'/w�t3_��)Y�N�/��~&�n�T���4T:�R���Nw�/@�C<	�������0���v�'�/�
�KJc3#�t\FS�^#��1���YQ��&��8{�21���v#�	��[ʛ���-� `ĉ��p<��/N2�ie'U�p�:��紙��Mei(0���Q�/U[N�6	|��S���nϦ*��ޅ�7���`��ph~�i{<�Ru%��q<��ڕ����ԟ�����u,�"8��>��4�5Ȫj���D�(�j��7��,� ��SK8i�4����)u$�es!#��4?�~�7'��l�u�fE��qOa9��y�[kr���I����������+רur1R�(�_���_j:����	�~{���F:ѳ�9^p��u
�5�Ͽ�Г!@ĥv���4g���SY����/��h�v(-JT��w���+Eq��I��1����I��Er�5h����#,pcT���?�MN�B�G���ZD=V͑S�s�{�nE_��D��`�U�/yю���^^�N��gR%ٖ�_�xF�ag�~VIP�*�Q���@��/��=�1y�=��Ǫ*j����ҭj�t<��?
�D?�Sߜ	ζ]C�3�F9Bp$���WG�u��IO����-1�@%�����M��b�hv5��ݩ�mCw��:�H�	r�􉦭���l�f��s�^w��֏���G,���Է{!�ρiځ+�6�+U�D� \;�:>��	��pO�n�/G�F�]��&~2:I}9��V�D]K1I���f�El7�g��F���
Ve�pAC��\���@�D.s��iK���Y�<��{������r��"��<���pln�����+�����ns�(}�Z��'�hQ-�{��ד�7�<��S��~~���(F|��?$N�*�g���T��ҩn���~��?,�����)�ݻ���Wd*WtS�"9���L��I��%���!��B�i��K������64�N�\R2��l�|6�S~$���x��K��ą�Y�]ͯ���t�:�x�I0���-�4-l�(��@�k��P�Ͷ�.Q�loJٌe�x��̀'b ْ�Lb��}���p�=v���!�w��J>3٣?w���M�{�'t��?��,F�'���)�_29��'?�؞����Tp�=�A���1����h�]8+zҒ�p&����{D-�q)�v0I�~4P�X�j�f۞s����Y�0{�HXO�h�ߨ!E��Y�I�118ۍ�C�z� b��إg��},�W���4��Ⱥ^�[���9�����`�@�I��X���.���n82�M#ZK������e��ʢ��/+iò�<H=�W�H{��/є���؞W��}]�:Їq���T�GQ���-�<�7��9���%�>�C�qݓEE�M<���X}y�W���?a��?�{���Tt�\t�,�D����A?��;�]��]�eHWy��bY�b�8�$���"י�:��K&{}��<b�� ��������	�[��ˈ�+���N�	�#f���N���U��
��K��6���95��Ǘ'������& i�j7&�(�#�Ru��~�'����	H	-E�*�VT��� �謃�Nt���Wiz䕍�$���Y�\���
����#�6�F���Xq��յ��|��4���=�HA�Ys�Ã� Q�߼�z�L��=x]	2���*hNE���|g,��g/hWȋ�Sj�&C���lտ����v�
��ډ��'w<�-(-9}M7,�Y�
eR��eWm�2����-���I����ʕ��@`��Z�Us�P�1*�h��&���H	��� A����ˊ�:-˥��J�	�`c9`r=O���	��Q���0��s;,Cs��Tn�ȹ�a�};�5��mW`䬧�ƓzO�-V��}!�n�3B��֜�9��W��Z��&k66���pR���%R�$���+u�S�<�};hB���Hu����x�e����,�uH
U�0������QoQ�el	��P�~�!��!�4�s�Z�6������!��.]��@�_�*E��D� F���2D�M�]J[��$w$��.�?ΰ��Hz�^��ײ�����(c.t��e,6�5mL&|%�D���$��̈́�,�Ȫ����V���N����M-b�vdL��R��9@#�<TL�#�g|�,�v��dv�X_�X Lp�|ꑒWs8�Q��a�;G�]��`�%�K�ɀ*|��q��^�n!(�f���\��%l�E|��6Իf5��x���z��r��:Hs�`��4x����O)ئ{O��XN�h)�{��u���Aĝo� Y-�Xy3���S���t«�=<YD/�������Us;����L/�2�����
HE��ÛG�}�9k��^1�r*m�+����N'ʛ�d��Ul�4���Y�#41"�4�k�9|.�TF!��H�1R�����t�D��!Ȇ�H{	�7�>rnc�P�C*qƜ���(]'�vmA'������)��~���y�f�|���lR�"��l��'{?DS#3~��0��S�1
(%ו&X�"�F�Y�
�|P%���]Su p�F͠G iT[���?vy��ft�"co�X,�mu�F��d4��3�U���~.Aђw���,�)�C�`�*�5���D���|�L:z�Rr�i98.h�����t=}�Z�_�@�����R�ە��+6�W=#��t��[f��jM!���� �GOƦ��&�e:M^���dd���� g��@B�E$�������,��|�{��./y�g.Q(<�Ї	�Pod�����	�'��e���bO(�O����D/���mLv�2[D�?��g)��Ti��4��;;)�mq^l��1)v�#��w31�H3�.U��XP����������}�� �{�>�ލ$���`�[π���$?o֕,��<P>�\ޤ4XH���7�~�X�7�/?�,�A�Y3�O�(j��y��^��zJ��2��S��M�3�S��8Ӄ�1Py-M8}�E����;:cuC�w��z�0��/T{��g(���t���y������9(��R�������[�Dd� V�aD��%�]�� ��*��ܐ�.M�_L���
FPn����3�PDB�.b��Ka�q�J�����_�X��{�1�NrY���P{���r��h�3މ�����[<�N�����ʾ
x7���p�����6�����K�k��_����Kv���5�j$��Wl����W��S���@����0FY8u9m�m>��|cv)��`2���S��NQ�bDg�2F��ԷGF6,��'V���k�2��#5&�Q�ޙj���'���'Y]sj\��.P�o�K�鿄),��2�`�7nU|ё�b��ĝ���Hsn�G�����HRKE��2�xې����Y
kX�.�0����H.�ds㭶*$
����	ל��H��_�Nl�B)�b��`�lu�����;��w�!�q>�݋t�| =��i��Л{MG{�,2����F�hun'p܉1�g�?�\�J�g�����-,7����%��5d̛k�kt����(���N�P���*�GtG�WМ����~
�<rY.cG5lf���z�ޗ~�m�Z��H\^�����[�+�$�h%�������7i�jaXF5E�&V�Ӎ-��d��e9җ���!�`���ň1=��(��
�����;�I�BŬ�r���\���:@�s�GB�e+������s!l
��A ����8+;Iߣ-�e�X��d`4|���	�M@�l�<�>�����X�s�j��z������"!��&$�[�(j�i\��K���s��15�pzu�7�K�pZi� L�X�I�a�.��iL�}:�W��1��3��S>���/gۗ���W�k�H~3�aý��&�����ߔI驶n��G"�=9���B�:}��_kQ.I��a�͐g������ŵL-��Ltwz�1��V�1����Of��A���޻wUҤ=���}u��e�+�;�b���w�fxI��
�2���|�Ał��u�T@l��������~��6!�Y��%�
�A���g^Qd�%�����-֛��)1��}��@:U�\�s!ޒw����<�����f�2E����v�C(�I�d�@�*M�Q��b��z�z���@f��'A�����ޔO߉����;��"�+G��&�<b�����z�uY0D���>�����\,׎y5�i�8��[�(]�W��Ư ڴnFc۩����bk�9�w��E~'Up��zߤ���f�cER Ǟ��c�.t�(�����;�u��+q�����<'6��c�����8�>-�;4#�6��Ǆb��?~��a�)jU���U�ۻk��9�s���=��X|�:��O��)� �o_�VU�\J�)���ץU�/x�4��9�S���I
:�3�����t�pzry��^��lp,v�.]?�D3>T~8���+�"���ڧ�غ���ÇŅ��{�&�y��~G�ݰ�"C��e��?]%
Օ�B �SO��2iݲ���Ȏ�	��8�s�ڌHn���?�X��8���ӿ�)6sB�jm�I��h� w[�o�g����'�F�,�\�����=r�%؟2U;Y���d��aޭω�hN��+^�7/r�����¤�Z	-\l+3��*�FxK����1O���I�7Tk`� �m^Qw���qvnQ$��a�H�Q���YxÂ�qx�}O}`$B�6mX�i
Uq�j��
��w�5��՜yK)�n�xC���Ji�ڛ=f��A��E�C�C�io���s�u���v�/�>�ķf8�q;��|Q��C�|��d]�����%n�d}�?��O����p)�O#�b�:]Ö9]#�6$��1,��Ke���M��z'��3����%�L{g�x���i7� ҫ�j��o�]"?6l�et,�^���왋�5������+���YU!v.O\��3>|U�yԂ�׻�������YqrR��mR���h�~��k�bĬ]���N��w4%k����?����n����&�9E:oLZu"������Mѽ1
�*I-gr�6+D$�߬��Ӓ�GW{(�z�K�ZE���) p��	�#���3p9�����\�#��,�0RY+������嶎I8y>��_��% D���yD��k8�4{�J�M��L�mh�5������!�O���|V�2���=���	��f�Y��'F�Sl.��/-X�F2�m���"Ś�r]b�j�Le_p�Mp�ԙ45��f�@Qb-�i�r�*�$�������b�f���US,��|���"�����ރ����
���S�;��k��.��I��*G?�v����ވ{\nX��� N����>e�Aۧm-��DWurS[���n�|��3�a�ӡê�\#�UE��}�����^u��0�E�����G���僑q'(Rĉ�~��8:��hCi�v��?nC]>��Þc��f��]A0����_����AQ�h__3�@�W��KX�.s�b�e��%9�8��ݩe�%=Wzhل�Z�v%i^t"-5�����dA�r	l���6B�?����q��$���Kԋ9�7��[4QC�zt�'���]�ia�0 ��_�eon����2�i��&��
p�����d�쮪���+�:�_Q�y��3��I�SD+�G��4�}�/l&��3��!fۧC$h?���M8�`x7p��[i�Q�)���>����$�\d���C��U�_���՜�W*5=��=�;ʔiQT`���h-��L�h��x;�>�W��	e�Zȶ���9�mx��%ݹǆ3�
�B+(9
���1�O�M�5�$�{�c�vo@ݤܺ���IZ��q®�0^Q��2Ϭ�4J������Q2���%YRt�t��=�W]�,Y�+aڎ��2�?1=�`\'�}m��Q|��K����7Έ_�d����o3L?F�U��x���u\�nN�
G߲Oi�^6a����_��m��N$�Lk�ht�$�Q����ҫQ8i�
a�2��8s�\y^��tW����ָ�<�Jp�<�w�	C�������a�k_��kM9ڛ�fI0��j��VN�:X�ޕo�F���2�Q�����>��#�oU��peV&q����L2������'��F�\%�X��7&8_Z�U�h��a�tFE3��MH)`�qƷ�j�a�!~~�~5����2�t�Y�.��ay���4J�ƞ��#6��	��{&�g����z��w�:�'�W�w�>D,�go�����"��d��"�yV�Ha���}�	\��&��2���%ػԱ<4?m��vZu������ؾ8ͨ�*������Q��@�c���teG�
��N����p5H�Y=���Xڢ9����s��ݘ̆��w�-�Q�Eg�Z؎��l�/5���w��(�j���0��'@����TȍQ��W����B�d�c�v8z!��I\�B��R�<�cT�p��8B��
A�oT�U{��qdR�Dc��=$��Qڙ�Z�N�Ч�����L}Lv=e�ۖ��OH�5���9���!&(Jd�L���7�q9W̄6�,�\��,!$���4���V��?�&(�z�V3�����-�\�я5�a,��=g[\ r��X�r��I���PU���q�\�/O6�����p�T@r����6}�w���ge�H	{S�� �q�0�t<j���ڸC��Ư)���?]�Qrʩ�8�%�앀
���"M������������=/�)�ɾI��-9B�1o�s�2��&��]��a���L9�����8Iְ@��5�;�$�r���[���(d�H��ĳ ,��CP����W ��,�:���O�xB��U�a�ϻ8"A�62y�,'����9�lߗ�6�j���L��z��)4��������EA/���N��66����BFc��JM�d�[g�o}o�_¢�y��f�6D�.��S�+_��옘;bΙ�Ob��]7��i�9�_�B�@{Ak/=�`bF^O��2��2tX�'z��`���nb��Vx��v�PFI�E`Ţ�\�D�}C(��G���HXh �Us��Zy3�]���I���q8Et��&;���=�p���k��ڠPhH>uz�O���<�����9��E�ʫV���lL�
%�0��Q�\k�\W���^$�%#�Bl�B�?��szy�6�@V-&��D4�锈�yl�y�m�h�a��N����C�j�w�5�Y�����J������|-xl�_yˀl�B�8՛��pC�-�̐/W��]���	O�t�d];c����ܡ�dS�Q ��w�;�6�O���(6����Y�+w�|f�X�^/��)�|!A����E������{�)�>��z,ه����=W�{��Q#���z�K��WDlX	�A.AS�$���h�ʪh6��b�n1^�����~D��Ȳ�3�iY�=�*J�kpt��8�p�ߓ�nE�m�0r�n��Lm�c���v����3"���,<�_��|�$�V�v�ׂ����7g�}]�#�^<U	PP�Ni��$���Sk�P�l�T~D���ԙs��=o֙w|�t�����CPܛ�`�]=�%C5�Gu���0�+M��u�����c_�Zf7�&��T=��r&��&��ث�
C��WAEc��C�~T�`W�>V�i��_�M"�_�}mZ��e
�%!���涔pZ0�3j]�OʲsYm���C��d��o�߅"�=@���'�T�ZElp��j�=*׈��4���r^�J�_О>�٨	T��۴�3R!�ޱ�|MMp����D����u�^�>h�Q-���iH�o�f������®#ua	�tQ��)�_�(�h*;�}d�ƩF2/ֺS6�6��Z\�����F�e&^�������EIBk���D>������M q͚�ؤ�d��\ϧ2ż5g���SX
�����X��*Usn^اL��h vnvc�}}!z�Y=�p�`�p%�DM9(�4>���%�_��u����q0���R.M��7�.+A�/�%K����5ع7ڇv��g�̼��<Q��ⰋD�>��J�[�MKA��ںJ���l`��f/ǎ:�wmf��E�m�%�V��*
�2�.��z�a�2��.5���jU E���ɂ�#�����;��ՍCs��~�Cp˰�_39=�,R&�њ�dt�NWBD�םR�1h�p&�����.Wz)A�N֦|k���ڲY ���[�(
�FT�j}����(�㰝�h*!���
Ma�w��{09�O1�x�^?����4`w �Q�_��ȉ�@��(P��Ӑ��gVV@���!�F{���'�}���~J�T���V�*����#R�i<Aw>�Fp�K��Q�I�O<�����rߢ~Ar���7��k=$���N�	,,����'	����%20Xq�)x(��8��3��p��9t�6��2��|�a8$�%��O�N�[-�m�6D�g#cJ��8�52���<vߜD(
���$.���<!`(��GPO�L��</wo�t���>8b��pi���NR���@�I�v��yKT�UR��q��	hL� ��8��'��p*�>P��Gu��Z��㋔�qʗcC�t�+��k�{U%��"�ZQ1����{=� ���� ��ә��}F��Km�?��}�.c�k��&Ը�TA �+�
��Z�g����?s�ȩ�K}�T(���j�"	��cv*Oɳ�>�		8��}NU5d��<Z�z�]>j������F�?��J� \.����Pڷ��*�)r翀L�C.>7��V05�fw� o�k��#�l�J\n�IZ��T�|��[*&u�6�7h�����h����(o�n)��&wS��h~�iyp�zu�^��C�h�:Ɵ�3MB ~�s]�zi*c�3@�Ii/g�g�� C�R�_���:t��ah����K+[(��*1 ��\u��g�!��P�;uS���}�e]n���*U��>G� v䆂�Ε�Q�1L��w�j��#�~��T��%Ć��,�}	<,�e?��\��@�L��860 �G�f�f~p��s�o����̫F���s�A[�*�5*�ȾQZ��'m�ө����W��:��\�zYg���;�Y��5&�M���H0�b�	��qqi� ��Y��!G���FP� 
|AB�؄����+�öI�uEr��`
����j����-�\�������?�;�/qص����'+�%w2��������ӳY툔H7tWy��g���J�� ���Â�	^�9��Ԏ��F˛�!s.�L�g�.aڤ�6;�<�u�E{�q����"��k��L%TQ�٩r��|���~JA�u*�?�카�^?��w�Ԁ�[�k�%'F{�#�7:b�{`X
��00�Kk�cI"T�4�CG>�
�!�?�a�ՒF4\��U���+DB�u�=�<����̨ۦ��bx�l`�%W7\�ř��Ț[ܲ��o@��} e�N�&���{�\	��	�m���:� umc�g6����-�4���}U@�����g�~ЗD�oP���'U��tW(�2ϔ[�uՏ=�QjᫎY�>qJ��\�Aȭje[́�l�w�8�tg5Q���|^��Tj'��#�߱K�Ph���Ϗ7��Ŕ �]�H'�fi�ʏ�#¨�\ܔW��kl�R�59�;T��.?v���#�e�ˎQ�~ ,}ϳ�_��X�`�-a7��w�X+�u��J�\����y�P��P|��0B_bJ8Wg��˞�НrF��7y
ǐ��?�P�?v��^(J�z�_���O��ڇ!�F�n��ZY�VԎ�j���t��qV$��ፆG�Z�J?E���J�Xut^1:��Q�	vM�UY^9�����?�0�����9�����#J�C;��\�Z��)U�k{�M�gy0{z���C��5������zq���0��U��}3S���bG�~�XZ��]T�K�������̮y��ǡ�f˼Az�ܰw�*����;]��A=�=��e�������J&
�X]��
ؤ_M)�|I�c� �,l���>
k� �	l���7���2���b 7¶A��p��ks��F�8?����,�� �b3�N����B�`Ai��U|��0�(;��8Q�鲌��$n��o	p�c�:x�V�on�C�ǿ�͹��O`���`��/�@;ٌ�gH�ՁwY�L�b"�������fOk��[$���Y%�٨Fk5�!�2u����i�E���9K��ɣ���Y(O��5q�1����i���b��7i_��v�/��N�z_����	зP�_��-�!����2HUz�#����nv����"O�_9'���@I�@��95Q:�:�o���A�DF�e:ib�����|b���M��PK��%�X�/0�\�q����BK�A� ��@i<D��zL�7U6�7�	�4Ol.�?&d�b�^E�4�XrE���<%u7_r#�j�n�f��2Q�.�x�ћ>���� ]c��x��rޒǷj��)	W��aG�94q$v�>H���*;��x��^Tr!��l�A?-�����W�-�v\E�������z	���9��F�jy�/��IO��Ú�,�=��(G��$�bw�m�/C��{�=��o�:���e��+C��-JSf⪅�H(��<�Dؘ�6�wwZ�Wt�XV7 ��dF=�}n�!�Oē�š���Kz@r�C �t ��9�Su¡RG�w�m�H�B*.m�xr�I���Z�re�Cb���ڙ^�;�s���*�� e@"_��o��+��!�)٧'����P��)-h�X��'��Ɏ/�Ҽ��c(�ܦ����ۉC� =ܷBj[j9�aT�T���h��et�>�+�l9*W�L�<�˛�C���& �?yt����%�pg˿ֳ]Yob�97��Z|�h���d�c��D��n�K�����q� ��; �;l��z���<Z�T�
�gF���#�ܔ��=�B`Fk��J��?d��#�7/�ͱP���r4�1n��C&<�A������a��F8s ѝ�f
Mi2T��-�B@�
�\�Ƚ��]=܊{Խ�r0j�(��+�J�l4���y PP�J��^��Ŝ�c�"�Y$4BO�y%WQ����)Ց='�ǜ�gWm�"uZd�	zn��ߋ�n� pЍ`����[r���A�����ZS;ݍ�б����lw+v}�(�mA#�OB>��l'Hiſu'{eY�6����?Ǯ��<ɧ��f�L���J<����@�-ľ�*���4�2�Z�4`Q�"�Gw ��`;X���6�V^��ZȽ|�/�4I|�/��m��	V�;HD�OWFt�����M%������*8N��k>�i���4n�q+���8Z�x�qƼԣ�ˇi��s`Vn���;�C�2iV��0���*����[�=ˀs�an���8��=��\k��X�׶ND���%��U@�^"����a)jq�H:۲ҡ��E߮�Sm���D�B���`VK\�̂���4ćdŰo���\���j�_��#ý�v̃n�bI���J����|*Gg���
5�ɢ1�)ߚ�?;7�@��ɎK����g�L�-)�{��3��yU���iԒ45�U���	�/��c`!�Ũ��qO�r�� �b�D����S�-X����=�k/w-�(c�d�'Y�=�,���㬝I�\��@|l8�����wK�}��{/qRz�AK�3 ���`�"X�y���eq�v��A~�{�Ӗ�cT�� �yA�l�V�m��x�~'�1E��BbTݞ�L�fU4w�]][J�/2��u��RZ��n�p�,�R�/�=YRۡ����SL0Ç ��'��|l�pdd~,mۡ+�7�����3�Me�������u�2V �oUPF_�lU�b6����� �ݯǅ���~7r��1���v�_e{���;�b�<m�.�[�`*�]��~xK���F�DdYY���쮨ڱ|'��������$�c��_� J�'Y���k��d����D��H��uT���^�9m����E�6���@z�lj�!`��6�n$��	��(��ʬ�5ܸu�w��\�d ��i�we��/+��J/�� �t��/7DYK��@��M�xR=���E���x��Q۳y\�j1M:�SΛ����&oDvpC���.������J31^�K���2��B���%�a�zKA?5�Gʉ�{�h=�=��B+!|>���<�ԃ9f��(�c���� �~� K!+��Z�O��s�/�W�Ӕ�`�H�^?�XS��� �ec�Sv��r��|����L�ȁ��	Σ�S��q�I�� )�e��S����sdC+(s�"�G��1���{�f��T`ؽs��h5��v�`mԵLp����ٔ06���Vf���;��l�Φ�_I=��"���(�wg�9���=*�ݘ��)�����/���}uZ�G��tt2�o�U%��X0LЧ�tPd ��&�d�% k��;���C�ȫ�?6!q�1������\R�?��<�������)�;"u�[���r#H�껇N{;��ܹ�0���AR���	4"��#F���R���{��؃��B�Lc����e�(?\T �@p�K��RYp�`6�5i*�Zgd�`��Ɋ�0pR�@�"��x�ʅU��(t8�[D�i!ːK�	�:=�9J�yW-�n�-�$Q�{��V�y�|�kN�5�a��S׹�r��d��Q�.u�T�����P9.��nµK����߿=	��8*�[?X�n�ऋ�"u�+�P�nbt�Xa�\ʻ���}@I=-������΁�Q�W��pVG?o����WZG�:���?J듫(�e�pد��d�fo�����^����^o��\��t��|�f�$�q}r]FC�]�Q=[0�	q��P��P}gW�q�]�X��f�����A4�U�̻=��g(�1N���hz��m͋�q6h��`�i��Q��W4�����v$I����3W��뗌�|�C��~�6��X9�٘-��\1/��Q��t�~vGI�{�������^���Ԏe|@4	�<_�eS8���l���w�ωS�]w�?M���M�Y�	�/A��5Qt�T1�qĨN6]"/�_����� i�ʓ�<��M�b�a��bʻK*�t�����4V]�x�ڄ��K\S��e=�s��Tv(R?	�>�H��r�Fu#"�$�DE
�0"ao%��b�Cn�b�\yd�p����	;|�S-}g�s���/�$bO9����U��aQ�N�����8�\ci.J��f�y����
\5�??�g��eE��o��f������g��i|~f/�ai��Lo�m���]�5Lmnϲ�&�9Ȋ4����ʁ0�v�HmA ��'��8$*[#p�\���]���A����-�p_e�~�q8�ʽn�x��K�E[ ^+_����Kb�ӭ���/�6a5����]��2¬�-t�Ɍ�O���m�E�v���I� X*�!��� h�ܯ�|�r�%bl{��Ŀ{�.�T
K$͋�+%M����s��(/�F
�çགྷΚHPf��^��Jk��/T�2.՗�+N$�}Mp�,_=`pj�Z�y�g�G!��{�,�ﴶO���[�"^��ґJ��0�}#!5b�~[1)����w���l�7e>$���	���*��ۮ�s�r��i���T�w5��v3�Z��PջŠk�N\����R;�91ƻ~��|S�k��P�1�F�x	t��f,L�>�+0�Q4a�Tډ��x:&�M��~���Ix���E@��)�J3r�䕷��`���^n2�� Fd��R/��o��:B��qw�����2�l��ۿ��@�E�^˴����=�o@ m����g?�RN��(��4�(ؒf&��]����.�OJE�5����"�D���Ǹ ջ���EKh���փ���o��I�/{3�@��vY���0�����[V�l���z�M��x.��dB��d�]⵻�s��Ղ���(�j@D��6� nK���=�Ճ&��{	k��VP�f,"�[�F�+.ȡ��(sgN4l�.WyQ4�j�i!�(�H=�����'��������� [$���["���FӘ�\��"�?�,i�����Z�Ч�DU��p���kMtl}">H�L9K�9q^���?����X�u��h���\��a�����q�p2* ^Φ�9c0�7Dշ���* �����
�|�*��x�����C{�ࢤ )Ϫ�^��>'@{7�-f��[pIW��y�G�p�'�áI�k�-"�>�RqS �&5�f�yj3��́��yF(l[��^��t#�#�lh�Ju�k��G����>S+�eU�7G�@�#�D�����\;�*x�����҇��[$՚���!�A��ߡ���q�@�Lq�}��9o��\�f8�܇́��(]�#�,x��@f"�!�i���lҲw���c<Q�#�0+���)������ڪ)�����(X�>n�7J?�ߠd��6����O���$�m�H2l)n�}��:�aG|!Zپ�-��C���]s���_�,�Ad�|������#�t=��A񂾨�>׮8��$T�����҈��=��Nأ$Y�JQ�gx����&����A��_/��W�Օ?���Hg=�t��b	��V8'D<D��a5���=&�b�Rfq�[��:�x�o�������f�ͅ�P��{����x�]g۽t�.�7$?R��O�)7ڗ�s�)�b!Ը�)D�(`?��4�z���௧�v�^l��7�WRly|����g���n�Gh7���<���|?2+��y��i���@��.�`��J��]n�?>/&�S����D�p
g�n��0����"K(LeQ�ou�ٱ���Է��H�X�2i��>hq�I(�eg�Nܸ��ˠ��;�`$��-)��,t��-�f�a_SHC�߿��aֶ�F��xz��-!_�g�Tpƿ6a�=r�&�{ j�9z�_� ��� �:�T�-Z�=��C|o<����&Fm�'�!��l=��m�v�)�]�wi�O�ɝ�lI�b´�q��R{v�P�;/��E3�A���F��t�}���w�=`,R����0�0B^rh#0�NJ�<��w���"�#H�{U&nH}Q�G�3Ck�@� �i�{�pD6\��Yp��Q�!����]�ayLºE~�`���4�S���Xn�\����'�p�X�5����N*�����R��sO	�TN�D�&��<A��������\f|T���O�9�{:�5W�S8�J�������u�i���bv���� ��Gb�Ā�3E����k�=o��Q7��{��㸶�v+%$Oq� [�Ȏ9�}��1qF9��'vW]e�����R�{`�ՐƻJ��dC�����������	e���w��-�Q��AnUˌ�i�4H��^һ��l-�l�S�v��,�_E+0T�[��֕F򍨬�4����M��;���|'g��K(�$B��C�pYQ�TV��j(xQ���_P��8���Q[ܨ���.��'OI� ���t}M��͋���܋���Q/���*�{( �����B5(����#�2DS�+���=yɨ���Ί��=^�������Nm��1N%�)��[�.�k�("��RJ��		�cߝ�e�*{$��d#s�,��mo�9<��߂��5�&(	��b'<f;���V�gI��-RWU�D�;�zFF �Q��7N���2�?l�<���өPJ��ӹ1}ٱ{k;����Ec���5<��-�9�dy�|�a!�#(�|���m��Z����-!����@4$s%84Kn�P҄��Q��!��_������[<�/3⓴�������0Fs|�	�)���]'���;�u�zگ�6Y��<��YZ'����'�l�YR��Pka�H�wD��Х��쟈�I�1<m%H��[�_�_2��__I%�Ta6s�����M�x��D�k7n�N�ǒfG�p��@Ͼ�_e:vc��^�U��������}�Z�*���]X�- ��ԅ�����^�ֈ	� q���[�H�����y�	$����G�	�A�t��H%��k�P��4�mBa�*�9�|���j��li8��3���7 >[�z����@����Q(��i?�<��2�_�g;�vG�ˌ�ݴ����N_TA5���u{�+M�nt��[�>���f�C帗@���3��YG�[k���P�]����K��P^�ބ�B
��e�	ƴ�a��������cZ�M��`�X[�@���Au�eݽC�#2��_V���1��sB��Fe��Ϲ���I��C���5����2P��O�ao�q:��쫨��c7�I�Jx5�+��U�����Y�f�☙g�����r��FPA|���o�N�����A@��A�"�S@LM�HU��wM����7���#'P�=�.��<-��ڬ�B�cjf�p"��=H�Q�UfJ�2�k��ݝ���6Ԝg�~�)p]�uwU����e�-F�����} �Lqx�\���j���H��� u1?UVN�l��<0Q�\�\F�ү}��'�K.(FV��A���t�o�l�'$�F���x�
��7�'��QQ�G�#d[ʅH�_���X5
}m=H��b�>�&�`B�0���P��g����b�n�isf}g�!�t��}��A�R�JSg�S]y����o��oɥ��_Ԕ�����7�j�����4�����MaQ�@��U 	\r�>:KȈɶIOlo!n��
��~fT,j@����D�jS���*�+&#�bK�#��Y��sF�0���Aѓ#��1T>_��a����羐�n��N������R��ƾ�{���*����KE�Y�<��Mm��j�;�7�i^���a���	�0��%��Vq��{��Et��0[����oI���N�Oe���������5���?@�	��[m"`�]�YV�d��{��l�jK�k��m���퉫��E�λ�	T��$� d �w�Gk��PP�i���a�1�Q��~�Y��)�aqk$�d�ދ��S�P�9��o��"��`����"�j�Uڗ8d�%���=��r&5h�c�)JjT���WV$ҤH�p����A�踖��3����w������ߢ}���ؤ���V���E���
��(\z���t*^�C�z����F�+���k�v~���.=Xx�j���|�	���V�i������,����oLr\��+/�a�����\,�a��$OC�V!���#����%j��������R���ʢ�������2���w�5m�m��S�蹴�1_ӥc:��΀ɝD�H��K�T����Lt�� L�W
����S �������0�0x�Mw���Gz��}�|�iG�$����fM}�%>��ʭ�>/J��k��N���D���O#
	��ʦxΥ<$�"�xЯ���WtO��\ۇͮ����M��gդ%+J��i�4�o��ZF��Y���t��M�K['�5�_���bT��q��֐�J�HC=�ܞ|w�-�9��'��5�����hNA�5�k�gX?9bQ#��M���*V��,��P���'ߢ]��������g�ġ.�<y0�o���2�Oŋ�.�+ L�d��xl�#A5ݲvHU� �ƣ�V�ǠX����H�Gg�b31kI���V��P����K��!�� ��!��hv��(���b�ܨT�XD8�ˍ/���#Sm�iL���b.�^���౹x�ia��.&)�ha8P~���j���=�g�րdR:'�����0��6؍ӈ��ڧ�� t�h4/ż�>�@��ʪ�!g��o���m�J�U2#�r�R� ��͉�g��O"F�[.��9��s�=�?�%�C���x�±��Ol��Ȝ�lt"�U�����q�0͐=���z%��KP�x�M�7�:S���G�j)����M�z���Fs��OKV��`�1p'�z(�E	�9ê�wL���)�_��V��n�.k¢h�2)���ÌsO̥Pw�L�>�g�8�h9� \$q�pzgy�슶_d��mẖy��$9��`E�9+"}>=�Cq,-�P]?D��qJ�+��R���x r~ܹN��;Еo9�"��t$*v�
��gU�q�R����� zSwQ�q�?��g��èU1��K̜E��	��F�t&)O����ݑR<�Rb͓4��_@�P�v0�%����o���7Eh���[ž�`X�F �8���1c�_ĺ�W��#����l����P2������������[�PG=��X��/��R�i�� a19k���B�L����@O��<*�s�K{�'�S9J͏��q=����?Y7��nJ�s9�\^@iJe��� _���2Ϸߜ	 S���s���~����A�q�z��K��(4�^�fyN���
VXĶ�� N���O� �ƾ@�e����18�q��?g P~dkTЪ=�geE���lN`���F	�}Ye0l�y�#Y][��{H�I�d
d�c�x�c	������$��������^�/��Aٕ�RH��d\�È���I���9�.�	|
X����+�d�������,�$���]!/��!���GM��j�,�C�>' �{VW���N�F�p��f�(�ᵿ��P3�Z��mk�p���{R���l�Q9*r=e�����dIwD�K�����H�Z#H:�0�tj���C6��+dZ��Vx��?���yn��`�e�0������4Rj�����c��ʭt9�1k�������7GߎW�!�O�(G.@�b\r�J��vf��H y��;���u-�6��y��KCixe銗o��,�6�-�@�!��~���Z�m��X�{�4 ,��y@���,;���^{��9�*?ʻ�3A�KY�M�BA��@M�ɕ��B胆byU��G�<�eEץe`����,��T��r��xt���e�ci
?3WP�RBRD�6�#��tNmuc��A��(�Б7�(�����P����5���&�n�L�\���Fʳ��\'*��IЃ�mG�帎�w�px/��9-v>�=�5. A�pu����b2�(Q����4��A��A��5�lk�n��������tHAO]�2|�����w��"���� 뗫J:��[�e��c��t��r/A�qJT�ݰPC�ߤݭ� +�8ްe��Z�K\-��dT+��	����i�6�k[�����a�wt�|�rHyȏa�'~6#�}�X��n���L�$]��*�>�r��9:�ּ��H7w1j��Ш�О���$q��[˫��w	���w|��:��py���	(� |;�K�ky��>���Ń�W$�e�ΉI�b{��J�$*���+�T�	~��`<�*~"5p��9 �
%$�"@vÅ�t��z}�:�Yc�r�<�0��s�����+ s(ſ5�Y���0���D���	T��&�xk:�	���<"��O�+j���Z�� ~��阠.3M��x�9�Hᛅ�Sw�`��n�mv,�Das�Ǌx�U�Ej��s͏܅�g�\�R�~>GL�4T��\�H:ӫw9�[1��;��0��լ�G3�_ɸGC�W��Yã/�iܜր���tU��&Q����U�=FP���;GdE@�w{�}�+
��r�L��!#h��YW*�i��Wu8�i�ˮ7��I��z�x�	^�{ZJ��U��E_�^���jm�š���e�R��"�-wKl<K?.�l?l�,1d񫰡��o�teK�bw�T*��bXr?栻!���di�C�Xk?�}>\�]�IK��]'�\X�T�2,�$���E:���&��r5R!n�Exh���fp%�:ы��P#{0�F�}@��i��seM����+E��
��<6�������������A"�2ɢ�z�o�rʮ�ߛ%�7�人��m� ���"$$KA�9A��SѰ�^�V�F˜�Kw���ɰkݩ���\�!9}��;ω�&5���X��\��Aq��)�Z�Ir����L�=�^��<�	 ߱� .��Q}ر���p�ּ����S5C�ą0���~of���l���mn�8k^D`�?bn�S��	�����\#޷����u���8R[��͠�	��D�j���Y
juj+bז�f�����\\<��	��ԩ���4 ��^�0���?��'+�՟[亣�I�G/��d;q��>N��Y�)�L�45|��i����(N�ٛ���wЙf%�N��;�An#)
�:M_�߮���3�)�y[q��>F�[f�U(C%==�NNUH0w��)�N�}�����><����Dc��	���-�;I�bJ ���L=�'�Ä?���R4˽G��L��.��������+ǛQ��t��Ě�����\T�G�=$c��O���ӣG6���6`��n������5N���6�Z2�Z�o��3�6�2B�TI�;r<�0ΉE�Ž��b)�!��X��3G�쉾�I1�̱��C��C4�$6�$�n�pU��u�� 4�(���������d�����c��$j�:���� ��w���!KeP��+,�U��X4��<�r.�.��G��.Y�Lժ���������7�I	3�oȝ6��gr��큪�|>��ɷ��M	���{�^�O���j�I����d�f�z�H�1�R˫����zK%�`���i��X��]�?ea
J�q2��]�s��7#uY껽驀򙻵tu����	�Vՙ���cm'KPuQ��κ%�C�=X������f֛n��Òe�%����6OL"�&��(���5列��i�gل���R����+_
Gn��ʛ/��H���.�S�:Bc�/I�o$��'_���6��m'�4G��,=I�=���W;͡἗U)2��9�/ݝϟ�̏��Eq�9�]���8�=٢��c����kUVa����g��� iN�t�p��ƪ��Z����'k�	P�����`�l4	�`(6�`��j�A��)�0OC	)UNE��T_]jU�.������Ip!�C�����h��{����X{Uw ��������B��.:���W�Xv]�.Y��Tu!�����`�t��'�Ο1P����A2�o�Ά�8uX>��$X��sܩ�-NC;a�]�����ϩ*��-��}^���<�g:�i��|ݰ�s/��	Ug��8����~1_3������ÓV�r ���fj{	-K��ܪ~�����9d�'�ܛ�m�˶W�&�!�P��'�R�&·;nÿ�q/+c��tjY$oRHU�m���G�?0���Yp?EO\V����M��@)�5�<L(���t�3�.v\�9�C�����m��{a����p�Β`���R��E������gK�:ʪ�����}U��T�F��;�ݍˀ�T5�S��c��Z��DS(�P{ wߝփ%���иt6�S�
���X�\\����J�)z<������d�vg���Ot��W����Jf)���&�5cV�h�=Е{{㗳�7�/ckik�o�U�ŧ��-��aV��CTͽ�QHF3����K䏍x6����0�BO�	�`3�%^�ݜ���bԔ�kt�~$�vN�䁰3��Z���9�L":��J��񪝛B?��]�`����_#�XbEcN�B�B�`
�\[��?��& ~[��8��hP|��{���o�f�1��ZQ���AW��u������%Ϲui2m6F(cGy�X��P#{�g��Ѫ�i`%v�Ґ��_�D8�7��В5��Aħ;̶Ƿ<�fi��j�ɩ�`�v~+��`Ps�'�IH�2a?�:}�_�\\��zR�}���T�]��M?Q4П�>��X�o�n'�;�ca�o���klUb��b��N�'sah�)�`��Gc�1����gJw;9n� ��|��; �cb[J0p��d�`~�v��}�	�s˕��:ݮ����o� e�n8�;�E���h+�2^�� G	��	�9J��L�8-����� u7���JXД̭1:ntRВm�#9��P�����$b���^��/t�Cr�[#3A[������MX%AuU�ܘ�b)�KC_]�R��!�!ys�Q���l@���D�h(���v���N�V�+�.�n>���,�>���!��mW�֙�r�%H�7�2��u�%�t4AUR���H�l��	�E��������dY�C���wVWxnD��G�L�v�sS��<��:j�	 �6�:$"�����{�X|��;:@�3�+M;��At?9���Ev��f�CY�h {�����ccG�޾����ܠ�
$I��W��+5M�P�ϩ�Ը��ü��wS�'/�����}v�5\k����n�Ǝ�(�HͿ�ףBE�Ww#�]���2��B4B# ��)�Ȓ{l�X����%�7|ucب�з5�g�S��MΫO��7�>0�_� �\�(����]�"[[,�CCf�����#a"!~�ĵ�xk�r���W�:��7�eԝ�W�^�s�`�p����YqZ[�Ok����ڭ8�Z�~���?D��������iv,�14u^�3J��;�W����w݀C�;���H���c����]��a�1�AK�y���9�fy�^d�ς�<��m+����Ю� #7\4�ds��|���~��O�dU.���ǃN���{�]��P��
���7����ވg �ޚ`��F |���W��g��R5�ɋK3�[F"ވae�+�Z��`!1954d�bI�)���F��a���x^��=�)\�ԃ$�/�5�y����6ۖ�R(�������d�n�	�UBD�FAj���65������D/]<��_#����K��K	�
�F����GQK1����3iv2:	C��
7�����D�X����lG�c�q��>�ph��Ţ�� <�B�y��Nd�>2s�e��φrǪʥ7���9�<H��^V׹ἀ	�4� ��#qC+�ϯQ�B=��?����{��?H4Q��18���;�����ܣ@P�-�'hG���*�u�k�}�
��=�+@e\j;�>趔���^VF��s��CK�Q���J^��<�3����TN���F��d�t@ꂼ�?���24A���z0���� 	B '͖�r�ɇ�/ٶ�F��O�)��%�5��*	L�%�A���T��܍����`��h}BjC/�*�B�뀳c��(����Z{�f�1�z���49(��y�7<��,+���	����]�7̚��Ghzݓ�$IQ�vV�t��~i�˔+��h��V�Y�����^�l@�>�n��?� _EIL?҂�-��L�)����:4x���و�	?�m޽H��^o�xmlȩ���`8��D� ��BJ��V������a&zLG��)��rm��+ddg�U��A9��B�� oH��N���W���nl\d�4y_�K%�d֜������!
w��i�u��4=~�w��CEȍ��)v@�ն쉪>�]�&˖n��[@u�f���
�R9�J:'��r5�|!�>�u	��_F귝'�A|�4�D\�Ɏm3��E��و��{�_>��Q���|�k�^��(d\js��\vk�`���8�_o�D�FJ2�n��2��m�
G�fm��$�<���a6�2�o��3+�qQnĻ3c�텝g���e�CH��R�kx"�/R��`R[�
	���3�ҽEtqhԶ�pVC�� dȯ*�+�r�����C��V�.7n0��gD������EZ�a#bz�G��?�&F�K�x�p���$w��H���=Nܤ�-�.�A&xEL6���������o�����r��<j�ء��?1K`l�m�/g+jxymMI�G.F\m�"<����Y�����)�����f���7�B��� �?��1���&�g++��� ���L�se�jƵ�x���d��#�',���0��	�0��7aC<A��Rw���MJ��e|�;���s��L!��[WnA��o�� ��U��Op��`�!��1	-�ب����s����yYL���B|�����';\�=�B�\	?��::�b��S=�!�nң��S0���i��¸��)µ�I]=c��+e��g�5 �h׀�g�]�\r�����RU6'حՃ^��n5�6tU���jp�2�w8`��u=H�/���JVvȕ�{�O�v���C����:78�������<�֨&<Xk�1���^r��k��-
vK>��oH��*]7ʄG�u����>��-G��#��K�vp�Ŕ)t�jV	2Aճ�C �R���=��~5��-�aCA�~Laփ�;����P|ۘ̽6zxU�������(%�\�"��g��i���vj����ɜ���?����v�"g��>1�1�6⢓�6rW0f����'4�'�`�-�Y{��N���ZL(QuX�1�e�٬ �輷�H�I���/D=��?bq�$��س��Z��M���?[���{�K��<���Y�ՂT�~
�S�+�v!����� ���,���{o>7]Y<�i���[�U-MwCIӝ�%p;��o�� G���N��%������9 ʴ]5�nv"O���	��'X�`)+}�="�	B=�^���ڣ{x
��R����X�qD���5��P��:�(���Pe����β�Ck��<#��v�1���H��������=&W�-ĭY=H<��G2/s����Ӕ���|F���ۛ%4�-q��OS<�, Q�k~��ߪ2w|\�LU�Y�>�R�Cd|w�i��3���_��*=Z�$|@�O|�F�U��U��(����S��ԳrX��4}KD�6�i����%����U��7pj~)/��J���h~To����E�vC�(!�A!lw|��%�Tm�qY?�c�=�?5�l�	��7�R��	|?�=G:U�G�������'ş��@�IL$_+"��邾P4l�|T|2-�?�ȓm���㏲���}낋�oD-�/��q�L-�7���P2f�&+�Qy<���+�E�輼��Dx�v��|���Ȧ�o^-�����7,��72e.�0a#�k�H�1ʉ��I��'�N���uζ �Wg��4_א��/����E���Z�?RՎ 6EՆ���i�����PW7�#��%��|}i�*��װ]6+uP�eQ��ȺrZ�*�u'U���A9F,ϳ+X[P?ݲ�\�S��>K0��j����VI�5�u�����ș�ګ�z��Y+��t4�s�����}�����Cx��Cݰ���!�3_K'�;�h��D�M��"[z<<͙:e�#\r�Pߣ���}|2�3�_x/����g�e�k��jݧ���l��=yk�BP�g��1`��xA��fS�} ~�#��g���P��x��%����To�����xC�#� ��}���3��fp>`�r7��
�i��̰�S}{-cG^�����v���?{��%�;3?{1�_�O� �~��.�J�L��q��"7{��`{���XK!<�|��#���ӂEYy.���F?Jw��(��M��\0��u^=�����7��#�����10��f��a���#�vƑ-4iK����|����*��&�$�ͱ�6������K�B���,z�ҔFt�U��{gq�F�KtŦ����ǼA�\]��d�G�?������A����B�V._s�Jdo"‭�cY�n��s�s�|�O��*��}�mD�n�Hl"����T�W�I�U��Foh�)T`���=~.�J�f�_*��]FF�G��FU��*I@sDgJ���a+����A�Y�.��4zRR3���c憘ܮN��f�H�X�8L���h�8��L���Ɲ���E����D�Bj���!�a$f���tá\���$7.�*���_�kנ*"��� f��UA�)A�,�Q��;-����AL ��t��LxN�-E�{�/_�����u�����mΘjUw*_����g�h�n�����|�|� hU�Ҡ��X�܌b�?�r�s�y�M���Rv���%J�3X?�F�RgX&�t��a���yl����0�:��$�q���	,�	���H.���m5��H!9V.!p��2g�9�a] u)c�@CS������;�IҐ�.�o~&��Z�K6%K��#�Y��A�O�ב���	�;tj]�xmC���l���L�~_LѠa*��!���"ስ�iؐa��xEـ�i	�Dc��[Ȧ\��NH�W�'5�~�:���8�q*x9���S��)�u��+��mt��~��6�P��|����ڙ><��|����.�w�`GL���X���70W��Q�$������K�df�[)&͠��2"�r�y�$�ܳ�.����`�����!��A�	Y�v-�?�գD��y�0(�UH��	���4��E�����={|8�� ��YmOÙ��ȑ��*�1�;%Y~���� �r/B���,�����.$n׎ˁ�����9� ��zJ?�v��Y|��0|2�+�d�rKN'�+���f�_����(g�4���#1��R���*���|���,mTM(!�C�=�����+3ȒE�'���$._��B/��1sdQ��ꀱ��v�v��`�c�hBc�D�6\����ZzI�:(i}\�-�х�zb��8���B)L�T\B�����i-�eɵH�b}E/��WsO�����`hD�Z����ϟ��P�WR���c��S��0��r�n �������3��_ڰ)6������W���-sE�*O)���R2J[O �=�@e(;��!i;Ά�����-��X��\�K=�Ue�i�=��rDY��� =�'ؙvq�[���K���P4Ϟ,��c�@�;�鳡Hؘȣ�/V0�PZ�b��!^��@Z���3pm���B���Y�,}�DL�s�*�sͲ�����6�A�-]͕V�*�ȵ���l�����`����8���@?$�P�P��3�@�7p��[g{@����٤Z9B�T���J�Oq0u�:��bs�Z M#%v�Rqz��c�w����(I�0�G��l�0!Б�:La�z,�jL����K�=/d���!�k=�B6�D���F��hl�U��|p�?���e���N[�5ή����+h�
J��e�� A.N��b-��5��pA$C��i��MU�6�(�L49�u�"-����ӵ�Y���;ʇ��t��Rܖ�f��J�η����y���Y��Q6��D�W��	�4���BҲ5i�PL�6D�	�]qk�ӍC� [ u&Ё�f�j?(I]�l0�H,���ĔHd�-��Jc4 U�a�:6Y�\����?\Ҧ~��̑���]�Xu�d�9��>U�v��A8&��P��b�TCD�;�\��4��t}���i=�*����
�YuF+��.�\�|Hw0�`'%�I/���]>�����>`\)f%w��CE���Gh蓩{�ť�|
��N(���q�
�3�F�F��9��2�����b�#�������.���n�O����1̒�\s��T�>��a0Un�[�t̷�z�=�*�e'�;H����}���.������y!~����	D��U�.'�6١�W5�T����'8�}BrÉ:~r��*9��k!�������d�&:�I_4�X7�gyA�3���CS�J���
'�)���'�t��<��Iv
��B;����.@���ߊ F�H�|�J+���]����3)/ki��p|)4�HևTd���������|C �#�O5�Y��i�S/MC��,�i���$��+���\*��� �=��FO�|DJ���r���w���-��W�]���Cر����uK U��c��\�$RI@���-G�J9��<����>����d�osm?�$X4�)�v'�w���ۚ����V���E{|�ə!~��{����eV.��c㐣k��RL�[���Xם�>�]��]�n�W�P�����ķ_�b���h�E�s�r;4�
a�c�Ū�eB&n�6���S�S\2�+�HAp���P�x�g����T�l��Ѩ�J��FàY;�T��'1��0<.��c��ݧ��	0��V.e܆��=�^V��|b)"�R-h�ߑ�V���p�>q��~B���*����%E1��B��s��ߪ-���G*�_���ȼdP��E�S/X���%�R�$DF)�x��X@ݗ-�@>\��1�����TJ<"�d��^�RX�����L�� �L��P��9�	\2BeƷ��$�r�����aiŽ�x�)D��q��$KO,��'��ݓ��"�(-�q���W���#e4E���3�L��:}-.W8I�`d��8��D���2A6f�DC(�
c�)��#�.����RJ󀟷3=���ܚ7��Ш����O�m�p�a\w�A?���Jץk���j�SYM�	���[,�11������ji��Zה)�	�`�>v��,[���'qr��3�L�_��Q#�(F�I�f�N�붴o1�L�F��"
�3�b%"�Գ��(�͈W"��}hBܽL�x7��	J�\��Ed���(�����P�O�}������چ"���$�!����%D�;d*�<��*"g��3$� �� �|hZ��)���rk�A���TYj8O 2BcO��m����]0��>C�-F��h訩'����f*��0B��!^I��O��`Y>�f0a��憊H�Ka�5wc3�u��gB㉦�/\�N��~�t�P��u���"�yDI�tl�U'�������}&�f��� v���'�P�<uW͸  *e���	�����2��'�@�������|Ef���R���I��L��
�|f��Z�hQwC��V6Y�q�޴!�3�`�FA��g��<��M���z��X�ܠ�GMM�),Dy�$�!��\!��n�iU�,n~�`����ו/*3�H�\	Qj����/�����*�Xp�>�-ב�]�[[�4n��A���(�]r(�}_ �C������9�s�r�x-�F�5:^�/e�55{���o'٤Y5U�X`D9��Gb S������GtN��C���I�T�����B�N��-M���}��{#�N�Ve~����{q _D�����|�(WR���$�3M;���I��k��
sPdDoQ/�,�p#��/���r�����e��[t0�B�o
��M���r�^[ɘ������l�=1R�]�Y�&�iD��2$�C��$�<!o�+���0V-ܡ�����fJ����oak�&�6�19|ޅt�[�����,5�:��m�B+)�z/�5�^�#Nͼ�n	�,��[�iRi"�!�x��v������������~;�^��r��D}��c+��l�B?v/K�d����N����Q]������nC}�z)k%�;��#�W��T-�}+vLd,Pk��M<�����_��>&|���w��^H��Y�-ؒ�z�!�u��I�_l���'�U���rWV�W�J=YCբ_��e�L���cU\Ա�2Z贑&�/Q���Y��-Aak#!t�Ach�>��ۥ�xi��2����s�tK's�>��Fq��D"���Xc�3�p�^ꕳu��t-B�!>.7�i���2)�OÖf	ܖ�V�:`�	,I>T*8��K��5�?zXOwԯ��)�
�<�fD�,��?�$@^N��S�$�b`Ò�4Xd8����+���r����.��Dx�v�2&X���!��DU�N�!��#��g��rT����8�:����H�@�� �Y��V��c#�w�r����������QY]|oF�4��2��?pn��.n#K��B��$�d��܂ޞ'��BSX����:����fpqɻ{�*�B��A��tB�f�@S�[�� BI��͑Y<���MZO�'��7`��=9�:����o%R�[�H�w�G�i|��F��C��4�qH���\�=�OM�� ӌ�f<��o�}���)�yfl1��H�Yx
�J���훫N�T�D|/�q{�/�=z����tQK��q;�O������\W��cp�K���3ſ�ع�v������y$�vc��TK��G�m͇(�C��^�T9%���ね�Vrp����s^�I�C�~%+��L�9�0:�ed�]�5:1'�m����n2�*�"�`�
[����B����GZeE|�3-�q�� ǣZ�MV9w%�f��2�*�}!��T8r��הv9�R �$�E� �f�'ӵ��J�5��c����G�MC�lht5Q����D�K&4��}D���&�wtQ��E~�9�oe܋se����8��C�?�O$
��by�w����v!��V=d�4��1�-���ݦɄb��:%�����@�ɡ��%MDt<@{��	�7������)A�?,G�AU`�A+]�6�*y_V�,�����*���h>Ȣ<���K� VE������0y���v��W�@N@sx�����:��f�F�u�xW�ֺ��X��қ�,��)�J�s^��ĝ������i�7�i��e����?�(|���v�I������������)\��p��6���������o���v?�C��截~�g�k��
���a��Θ�c{�ks�xV`��x~Ϟy�Ҏ��ť.qLf�d�D����؅��fbz-�~CZm�aC�Q%� ��%R��OW�+/5�ʽ���c+��+,�w�	�J��o�@��+��u��*~B��ɖ��ɰ��[+�h�~*�����˲K2qiǱ{��v�b�tӈ]�V9ݰ���B����r���CB,!j�p)��T��.b�Z����\�z4��0J���U��Z3��}�4����$Ot�/E���O8V��a�1���B}�}6����9�Wĭ��zӖ�]h%t[��QK����
���-�m�>&u���"��<��7^EG�#�o�����z�Q��h��|%M���̼~���&�����gX������ؚ�z/K��8����)� ��R��.��ּ�,Q4��Ֆ#r揾��NK���̀2n:mn����MX��K���v�����4�f��+��WرkrM�5��M,��Q�9�4���o��uԁ;�*W����'!t�Uo�O��i���)���ʗ�i.�U���h=��=���!����Q��W4wҥ�/|Ƣ�~$~8�;y�T%]�zWK�u�[L�S��txdeӌy�azS7��XP$\]{T�pT�J�p�r�~ԗ?�Ю<�Vqb�����.�l&ߡgy9Z�p��B�{m�NFp� ȵn�����J3K����#ԟ���;�w�
��Cr�)��wB]5��Zu��/��U���{��УV��$��㙞�d���1 ����藌|�v�=�aV�ߙ�F�_xE$��]T���2U�D����hh�?��m	�z."�� o��Y,h�n���"�a�[�Qb�o�E��O��"�2;�3���_Vf�z?�@�zr�rWt�N�/w4��W2JzQ?��4̣���/���W�7��z�/��zB=�t
42e�^jGX�Xjh�/�����@���K�۩��Xka�V��:r0 �&� TrP�0��)�nd�~ �˛PO�/f��K����i���/���q��'Z�Lʏ11Գ]�T�oJJ��iYA7�}�I�0���6k3 ��J^ئ����jے~K)�^�,���	4��=����P	�V U���:ϧ�3@�?��&sݮMz�F__��G��*��bJ/��FOWڀ6΃�`�[���L���z��U���!LH���z���s����v��d?#�$3�C�����O��=���"������1
��yh?��r�[�8�r%#h��������`%��g!��ۑ��2�)7����/c�[��I���Ѡ�pF�3x��\g���c�q��5I�uޜ�@��
}74�
9I�`����V'[�5�`��;Y'yY2x ��Λس��{x��[<�,��'��"��5��(�����ꡦ5�68��'����ӛx ��a=�)�
�����v1��-[O	*>�W��u��G/����W�b��t����@����DQ�us��֦���YF����|a��ý:cb�@��?����tx���I�vqǺa���Ł���!`����M}���E(p`0S�����8Y�������E�|�(	p�e�J�ԷC���7�F{����9�A�q>�e� �jV�)�v���Cafё�ĳF�,z�L݈�t�D��Ҥ/�ݠ��#�tFA��@vG���E��¡ͳ�d��(�r�����4@�&sY��O`,#�>v��5�!�];���/��Z]��䇧�|N����;M�©n���OGD����I��%��$�l�tMP�N�����Z36��^�Ԯ�e��-8�60a@��m��㟌��N����sz\!;�(��?����$��ޭ����� ��.��K��H��c+`b%ҧ\�(�=!G�����U"�u��l@�\�sӿ�������T�HC'ǋ�a�䑍[v��ܖ8";kQ�.,�ձ�]XF��wG�V����3����論�rfr+�)�ĥ�W�0v���~�.@88�t�Sr�P�� (ԱuϘ�:�y�+
����*T�Ĩd�h�%	_�?۫�ߢyQ���/����w4�N®똭��n����@�*��6���c�!�|��nt��s�-�������)�&N�5�X���R��~�?)H�΁2�S��jDS�J�}��ͮ�i�t����v l8�*�Jc�2LM�$Ǖ_!�T�1�^��#� l�E�!�՗��PZ�� �G�� ��/Cz=w��b���S\�#���[ζ�h�
T�7w�Q�m�R�G��-f�Vߺ
L��}fëF�D��Z��RPĚ�w�#�09r���zݾ҉�����'d�ϋ2P�[��G�zzR�yqf�Ծ(`���@�\Q�����AI�џ�V:��q��%�iE�1�xom܅�	�Ȉ�ӀݲB���I��>�ض�L���8:�8��h��T|���Pݡöe�Y����:vMp:.K\�~���g�ـ���8�]��h�_^E�}�I�B}�fa��Y��f�Ԝ\�9p���f}`�8e<�w����Ή ��<g:e���먚����>Q����>GՍ��4d�{��}̘��^Vߗ.�� �4%F�p�t�.�^����<E��v�3�DhS�rR_zq)9~���y؞~&ndcށ\b�t�����:ˢR�-sne����s.� O�qN�y�Q6򚍊Δ)7�
O�~\��<��i�ד�u�t(ˍb���o���G�p�o�ZW)�,W�����u�A[3��l�#�P��۹��7MVr������w�ċ�!��n^�
�N��Ȯi��h�X2�މ�M�g'	c����PW-i�i�9��Y�߸����u}H��S�B6͘�m��q�+rZj�Z�i�5�_�o����j�#t��vS6I9g�$��D,��n(����[Y�,��)%�6�����3���	�qMj�F�H臵�Y�K�<d�K?�ދ�}̻���$Ac�[�� zߕ�� �j��Ě5R����M�$;?��ON�4���.��	���/��/�6MF�,�8�6S�;<F�����b��XL��z����#`0�U�7r����CD@s�u��3��V<��MbVlލ���X,!�Ѻ���r�bTv_m�
��0�
a�X�}�0�+�Q�?B'�yN2in�$��l�B��~d�{;�bL�7C�>�v�`䄜��,O^@3Z����n��C�0�@��ig�hM3��8#0��x�2�ɸ|�������~�r;�f}r��F$N~��N�PW�ڜNM�Mdݩ���zWV_W^�L���`g��qj��m�bfn��m�w�ī����y���O�K�_=�E2��}�Z�5d���Kq���2��:�����K���9p��Z
���U�]�Q�|�l������`Y���:ӣET�& y'I@<FnPj�X0�z�Gx�k�]�)Y���!��A�z���}�'-5�j@F<��ϫNS#7'U�r�À�:4�5\�KC��(��d�$�B`����)4d����j`��^Y(P��N�����H�>��3]Y�	H
~�-��g$�7���=n�J�+V��S�l _�O�ӌ��l�����"��UI��ߞ��������!V�w��6���&V$���Û�0�� o�;��tۙ;���i�lJ2�^��K$��n�KҌ��_A���'�4���p�`��XGn�!A"���ǥ�IJ3��+U����ַ�W���>�|W�r.r�d�5����l�"D�9�S#nZ�n>Uԣ���"}�K9LkM$�����Dk��\���]����B�?�7�Yٱd{!�ib~C��g'�9W0:��mO��v�`��Q�x9�l�/i��hK���ul���-����D�PZ��*��DÓ;�F*��ʱ.j#�����O�3��\��oL%�y�A�,��:���^R�rUj�d�z-�-A���t9]���أ�f��`�#���_k���f�{��2�7ɭB�cQ��whٯ�<zդ�����c"��l�>�E�,��E�mt�d�9̾���-�,/A��z׬UQ~��dj�rsd��!�K�:óGq �I`�����Fz�s`̒��E��7����k�P��1h1���[i�)ص�АX��yj�\Ol�i�S��9��@F�e	<���0Ǿs�� �tʵ�/�&М�I���ru-�J�#��d�Ã�Q�؎k�����UK4|,��Y���[-��������;���6,-�w&�x���r�> �{�c�R v���G�\�0�@R�T��O�o��I������G�d��� �vb�*��t���g��˃	#�Uצ% ��Y]Jw�|7X�u�׿O>�Uٚ�k1�|c��t��t��a,�EK���l�	�_og���e�#�P���)@QCc�p��JTV�U��5������E���G��k���e�QZ�u���λ����<lIH?�A5S>F{ �J��������I���e�Va��s:�4�ɗ��֓5x�|9T��k�I/��$u��5����397S��
�,1��=-�тG �iBÒ�2�Z=�#�9%5ck�A"��ި��y�?i�V���>g"}�����ya�/84�K[{y^S�5������a�$���p{/uB��/�]�6�cr?P����.P6X�~n�-k]�@+R�s�*�%��<���c�7��>vO�V�,o��$߃a��ŧ���9�z��K*��pG�q��b.ҷ��\%mc��Q���H�(9@�Аh�D�B��Q�(�AC�:�j�,���`�{�|��B'忹9�����Hq��)�ẳ|.���c`��Be�\��;��� ��H�����ЗH��F��֬Z����#��fLA����Lz�;��a��KrUϿy�Ɣ�1�}��
t��p��A�l:/�Ĝ����y�	�'=XDb����� ����j�֥���p�SE9+�ӂ��3���J7���P(IW�CQ�BH.h���񶾮Q@�YP�(�}�v#���P�lu򰁩 �F�4C�WG�3 [��oڹ����������>���ML���)_z1��}�/����@O�y��Ì,��c{�'IW\M����	]�Ƴ��f������2�yg��-�U/�l�\C�/��1h��k2�MP��-7vD�ʋg�k<�� 
I �MF>,�`8h��� �������v��p�{�$z"�o6U�*P�.E��Y���,	~IVQ��h�,넠 pwf�q�,�OX�`LV��F(�]�ON �\���b�&*��0Q��0�'��p��vy@�32�vP"��c vf�	(�(jf�آ�c�$���7��`�l���L�0*���)���&;�l��/����kc�����T�D� 4�	0����[Q�� ��!&_G�g"��񂾵���B"�Y4�I��b�p�H�aLcǒ�@;�0���r�/�"�i�0s�u�_^��<�꠼�s�7:�2�k��ϴ/p�0.�t�Xr$�q�����\Mx\f��\���h���.���>H�!��H�r���N��8��=�gЍ.k��fh���Ȏ�鼅P�%��?����6L���#!�t,s
��!�X���\[�O��(r���'B��Y��� �@��.x���-���H����j�¯�WGdp�/u��9�/N�e�Rlp�>�k#���&���?�>?���;��})�{��	ϲ�AmE̮N$6��4�~yr2s��K�n@�m����"Br����(�nx3�X���P/҇I�g{D<�����<�~-wo�#��2&JM�=ps�Y;�5�đ��	Vka&��̚U8Ԫ�:`|��J�A�^�H���L��E�A�> ��w��U�j퀕�nxch��l]���HF�I٦�:��=5����ˡ�ur�M��!�O@SZ{a�����˴�9cZ�P�w�w�t6~HL��"t����R���-ޓ@�������* ����PG;�F�f�V�����Ā,Y���ѱV���ₗ���1�P���#n'<�*��A}��RH��Oy�����0{�]2ജ��kX6�8��i�|�Yi|�^6�Q��s�e����ԊJ���f8���;<�﹊wl����ټ����ln���*�V�R:��I榒k-7��mʚ����+��^���t#W��w�4wКD��N{���=T��
�gn-���ca[`�zjYM�o�iO`����}!���kE@��EGIp)�Q��1�4��m���1x�a�|��L��7�~>n��"k���cE,1�H�q��N����;�2kn/��,�%��,���v}̕�w=N+ɠ��d-�4���6|̜����"��c)��?��5���oR6��h�]E���[��ډ����ͣ�<3]�A�Õ+lD���-�s���gY��F~��_�����b$$���?ǔW�0��x_Ԑ�?~� �l���1���y�O"�bu�������x8�m�f��i��8��Kݛ�=0�zw�㤚��V��v�ꆫ�e���Ѭd����S�U����"���2��s�3D�����I��i_Wax��-��ܙHB���KT��#�hԨ�UtV��-4��V#�A��VT�a����DTR�s3�Ɋ6��=���Л�ًV�@�[lE7s�?��و�}
�t(��
Dm-�ߪ:��`���-U��ѷ�#d'��]8�CY�FH}���|�u���a�`yYx�l�4e�\�"$��OW��s!gxR��g��d|�c	2���Ⱦ �@�RK�)�x��r�⍅oܡ�a��7J<��@��B�(���.�Ь�BF�s��d%p���{i�4;���s$��d����z��$����8˛���!<J�!��n����z,���Uk�t��Ґ�\����7	��%�b�5�Pq�5Y6���%�u�v���.-��9�kev��m��O2���p��U)e�4�$@:aWD�g��_�rI�FU�J�$��-y���+�����Ў,g��ٿ��3H��*^��UU�(�W�������� {*�7�6�W&��S%1��$/[��C�	��#A�Ib�*6u@ܢ1f�{�lQ@O	�!!T���?/�y��W[�c�Z��^fω�.�CV͝83%Z�V'l�9U�`E5�XO�w/�c�� 3��zx�4v{�ˈ�(r�K�(��iV<i���;^�� �w|�fA��O�jyx���n_���Rvg�fl)W�>�"J�0�WD
��'x�W
�I�'�Bx�����6l�PN��Ep5`]ɞ=�\��M�)Գ��#�Cz�Y����7#����!�ʏ0v�W?�"u|L;��QR�xs7`{��j�V��S}�h$��Q����NW�ԧ����'�n���f�j95�t���t(9`�+S����aug�#p�
m�H��.N��|���>5�?�T�D���Qx��4,���.�'`?���]�	L�1R*?����M4����ȧs9c'ui#Y?%�3�[7��\s0��n�k����tlИ��B�i�:9n���=",�A���Ȳ��B��ơ�>�[=�'�>���q�
P��+��)'�[}-d���`M9*r(��2(�Q���` ���<���SF�.�Lӏ��7q�g�:�!��%vS����ΤT���^kci���Jr���ÛKc�"�ŨnȖ������9a�Th�2���>�I�%"t�0T�YVhRڔ]ٺ�-N=�<���T�+;�^�pa�i	�Y�"�>S�}�3t�O��SE䀧/n��6ӫ1�C�C��ݐ̵QJ�g3�*��9뜅��c���:aX�j+�>�v'���g2� ��ֹ�|���M�J�p7����zD(V�D��lh�YS�ǡ|f�������,�]�]̈́Tj��b��������6�'6h(O]hqq���+&���/�YB'�2���f�_m�>�F�, ]Rt/������7��A@�4�o�;{l>�7!��8]���*�����-VZ�]M���Pn#=��lb��g�DU��24.��uƟ/�ޠ2�A������<�� l�y<�
vߑ��zʔ���O� ����9xy\m��Ƨi��/t�D_�֬`ܝu�+"����: E�#���&�?���xp���(����qv�Z�pP��shU\�o9�h%��*�("������HZ������ř��Jғ�+8�x�QD"��a�M��.h�g�I��I��jn����Té��)q���͖8no2�X^f��Zq� �BG��ߎ<thjM�I|�s���`��ܲ	�����W�ϲ�g7*cv)�J e��ͳ�㪁P����R����yr4<5�eE5�:ʶ�F%�Hf'�a�_]*Y�|�oz	��Q�KWѥ\��g��sb���"�w"�׈�g��6:�C�8 .���I�_
�]��h�iuH~�ae��A2D$c�e���5� |�pO.
-}+����W	R�z���\�r�Dj �h����t �ށ�ؽD[ږ�Fc&�y.!���1X�3F�xR�����0y��l�?�:ͫh����ǁ[Ȅ�9
�Է6���,�"����e��9?�����^�F��u7�ԗ����$��_f���=��S��F}��M	�,�\�3K�T9�v���Lk_堓���aP����E8��P��=�	��+��P��S��g+���U�����6FR�o{���k�[�_��L<K�!֬.���1��R=��#7�$S>�wŭ��w	�ς5�Uc��ߒ�zDy�0E[Ѹ=�n2wdK������+iDa�%ތ^�;wI�G'��5���]����ժ��Q�dT6ct����F�`o
��vwS�Ivv�!8Pv�&�?(׵
\�%h�B�G�ȡSwm�O/-a�!��ME�,Vm.0��d]�~��X��q���UZ�dL���nj�+�~.�9��eqw��ny~H#֯��n���\h�=-N����X���~v�u��}]`���G�%p)]i7����t9E��$h�\cֻ72V���*w}��!ʁEVtk��R�dt�:�m�1�7��sڲ�ƕ��� e�h�����BG�l3y�Qߌ�Z���6g��9W�X:��7����%�nZ�^ʵ��-���$02�βߊ�A8�p�Ik�7,�n��Ѥq3ʦ[ �ny��V��azwf�gl6A����a�/���x
�īZ_k�A8)�LU�Ck'B��E�ʱ��7��-�:�@+r�����pz20�NMBr(r� �\jX!�rT�����G>q4{nڇ����4M&�� ��]M1���L��('AP	i��t[Au���%���x�u�0|?����&�T�o49����Gs���D�w������Oℵ��H����㴁q�#��E���Կ�v
�C�X�eW�P��!b2�oz|jU"�t����/��T�Y��L*P�D܉{�ծ%T+�tU�l�Q����A����ari�A��˂�<��Ϟ��*��r��?�*��Y1�k�sG�:�R�m"%f�`�
����1� �LNJ���,�������f�6K9�Em4�B>�rN���;w�t����75Q�����N+:\��ڹ�{Iw�"�a����,g�́�	l��|	:��_�O��pg�����<�c8!�j�����Eg����H!�BK�H�pV����3J(-�j�ԡ��s\Zos��3����[>.gB�G��gUa�ֻ�Ƅ)3Z���������a��6c3 T:�� ��&�1+��5;��eѶ�C��6�^֘�;�'J������\�D��?7!�圷�($:������w.�PL� d����ʹs�"��ή���K�
.zS*���ǴY�r�Q^�D9Mr+2gj��P_
�����tL	�7�I��;��������/MO�����v������\��y�E���O���F���(y�.`OGbO!{1������>�gn�n�Z/��;�!p!{�*K� v�9lne�rBA�p��X���#��CQ$�������3���P1~���s�? �Ą��/����X�� ���d$0�2,�2���D�K�-���n-�%�x}�U�)��T{��d��In��68 1m���� 9�OJ��uO��y!�};t&,POt<��Z����!B���be���nph��K8ٲ��ϒ�/M^���F��z0��SWމ���Fm�B�Y�S�a�N�����Q��]��J5��pl\�!��?�&h�p�k��kH�rYv�����#`H9@<�$�S��0'I���an(��ؤscP�ӾﭪT�!��� W�FPjRp�
(�]����iR�C�p}�Uc��N��ݩY.�8r˪�G!��@7�c�G�1T�'!%y,j�ր��z�ɝ�!�t5Ο���(}N�|�p;�r�W��h���~���1�/F���U^�����a���v[ğ?��iu���I��Z�&�as�2����)#Y�;�)��d5��Y�ex�]�d쀘I��I��Z��ݻ�~��b�$~��YEQ`K�׿=��n����qL�X�Y���>!d����9��@~>�)����v%wC�l}f��Z�#�f!���ȋkZ�I�6b]\�+ ��<s�-Ap h�)���!�M�:��H�	�E��ߔ5�R.Y���rB۩�\�م#Yն��~���#�p$-*R:V�>�:���.w�;����x�w������XU���k_G�����r6T1�"a��n]��d��V1F�#@�nN�j�MJ����O�u8�<��8H�}�����w)h�|����WH��ޔ�pĩ��:��eѓ]����k�GL���O@�W3ъ���Ä�K�L���y���+�.�v�e�J̣�m�0�SF?��
��������#<�o�OYOg�6����v\��0{�2CY2Ė�r;4�D[ 9d��匁���i���0�T��࿎+���Zf�=���V�ķ2����)��q����=h��$�)���d�&�y�솟QT�`Ӳ�w%�;j&CL�*ʷ�e�\�(�b�jt0��i���Y��t���w;-S/�� `�8�����m>���%?���U�E��~w����@��t�jmuc�"m�����8�r�����3tR���1��/� �je��$�`!兼�9,�3`�Zʛ����>Oj�׋[��o���(�E��
;��ޤ�s����oDB�ޥd��xK�T�;��Za~\�|�E�_H\M���aQ��y�:D$88�V��yh�Tk��l8h � Z�z"�֧��� _��ꁱ$���h������y��Yx��
�� ��`�3�b���S�C�( �Zfml��&
J�/�Ƚk��_Nx��Xսt:��U.a�y����'��/�l�|ǑCl~<4���n"�����<��^.(�{��7�yj��J+|wB��f��Gq�{�ST�S�����ך�e�� p?ٽ��t�Sf�ӣ�2�u�:"�:��C�`BvJWA�p��~�d_A7���`�܂˰B��o�D@�%�U�ȗ��XC���k��}�������(kw<M���#z�[,ӈ�S��"��O�_���_E5��b�1��C���>��3\���:;��u����h����L���jcf���r��nۚ��lszE����fLШ ���Ku�{7>`
����A�*#��cƁ�`��Γ��ޤD�A;ݩ��|���~��)��A�A2�ۑ����4��[Z()Zz��C_��e��\�*�]�qtQ�}-T�58ULȰ��f^� Yt�F3���b��^Թ���#�q� =	��o�k�:�ո��.S(��D{�e:��Ӄ,�|�:�ŷ���O+��f�-��仓g����s����|�H���`훁/M.�,	���h�i5
S��ࠃi��5Rև�Ӏ���x�hm��}��#MgRm�o�\)����R8�s�jse�<��9�_��	�i6�{�g��+�����'�ٌP �]��B�R-ta��z��hC#�vhWT0��b ��؝�A���솶��/�
�s��[�a\ίj�X�oG��������r����	U�[����q��=ծ-���#��A)�J�0^tp��J�PQx©Qί�t��r��+>�Y�Te%����n8�l���BL��K�?�8�h���Q��
�d*w�b�J�z�P+��X_�/�\!Q7�/��g�}V�vԜ�&͆xR�9�ȉjxXY�"�����-a�$w*��`#\���r��i>�p��9�6�u��b�"�
-�!�H_���'g�Y�v*�~� ��g�N@9�e/�M�G��z��l���;t�é��W�Nr�
�ϤB �A��7�6��6g�;��S�'lC&�����$�	PCNʚk�SQ����zl�[>&,�k6y�v�6F�']�j�L�N�I�
�vWb�=&�L�c��'�S�!��� 7��q^=J�Wv_}@�@��������&qEbHn����~�ԳX\�[�s�� �Χ.u3t>n��	��2���O���S�1�������7�7Y��
m���#�V��g���q���~@��[���^X֞qGSP8\��Rc���7Qk-� ��j�8�ف��4V��!�~�Lx�^q26���i�w8}m`�&���Ip���"P����r�a.X��'tC; �^��yϮ{
،�9��V,�TͺIh�������bmk��=�����.�0[5>��	��W��Tڗ�@�%{&g�����T?Wd����4M�i�>��m�����vt�"&���R��I�!:����T�4�4K_7��^�L���q�xӵ��|wT��lIM��6A������9�cP/����1-o����S���\�3f�^q����qz�;����zn�jǵ\=������\Mȶ;^:�R�J����.��*ֈi]ُ�;B&�<����2���Y������u�k�t��AFg��J����k�g�x��1���ï�'������}ux����4��eSv&������<�.~���}�����Ut�� c-uD�L�[&�������x�j�Ƚ���tu�#���Tr
������ݚÞ������d���oL���,GB,͏�Ǵ��v���]��ts=�f�}�V}+���e>�y�� �-@���`��P��:ց\�#ı�2��q���F����S���G�.�}0[�����d~6v5ޕ,��/\$cw�M�K`���G��MCT=�`k�ٺ�Y�G#�1څ�A�щ-,��U:PS�4*�[|�Q��D�{��n�b��Ҧ���1vN����n�m���`Q��g�6v�JtqW�T@h��A��,^絮ء2�/�|�B��(�����-9��f�fY�v���*��"$\��F�>u'�qbY�u�M����5u&���W����~��}��V��[�(�4�r���?�^ga��9�=х��a3�)9`n����禳�ʡMK�Nzh�ۮ.��~�`(ₓ�0ߢ'��ߡ� Ӿj{d�|�^��%6�"Ž���s�/2):�f�K5��
�Q�E�� o��.�˛�tG�����${����D&��w��`L78���I$d�����[�RN�ջ��i #2"�5��Џt��(����x��O�j�I���
 ��.��`v�H� v7��J��I�ȡp�b#;�-0"`�x�~���<�^�-�(�\j��m��d�/���B"�iFrTi]
�-hhY��s�$�Cy4��|�;�}*Sz=[X����LuE�d����~�A��@���ԁ�O���̋��t���_ܒ���G��|�H�]���m��wQG"-�]�2'��p�qxY�	�9ot8�p	n:�Zh���|V����]}ˡ�RŔ���K�K��\ ���,��C0+�Kc�آBz#�T|�(A���;|,A3x���:�v�8�!���/�w�J�R҆��w9�Ǐ��4HLxe�Ră�l4qt4�F�ph��/̂�O�OQ9�'�1U�IU��й��Jjǅ�)�H�Q�y����ll���=�S%�1r_G � ��[���-l��#*?�C��<����Q:�bNr��^�VYK��-�ej=�����ߠSu���E�瞓+?���6�9C�蟒��h~��G�� �է��Us������uY.x��K̄ӧ���0:&���~�4z�x�/�ʛ$��w;�(�0P+�M��=�7�%����	�BU#��AB�sR|�M��d����֮����~ӧ�"?K�zH�%o�A�;^��)UL�6 �-�m�hن�98��^�R
���^�k���%46��)�ѣ~�p���Q�Y�>��5�(�'J��xZO&��!��2+���ZoW$;����������B�"QY�k�mS|u��&=�Z�jF�.�黢=��l�� D)�a��8z��F/#J?E�i��$G9M-��w���@;��|�1 Fg��|���՝�R��^�+-�x/2����dr���ю<�t���졠8�����E6~YK��F�i>�E�ow)bP)q@s� v�#��7��|<�����!�0l�B�/�e\�4��RP,����f�n(>Q�%e�5.��\��D.�������0��ʜ�'��ޮ~���0э�3��|Ĕ�且 L��$˂���z�]���D�cK���f�2����3g�S���s���4W�]��cE#{���F/�~s�\��8���l �g�~ۃ�G_��Q�}�`���@����s,ebjv�k���c@kT�9*4�.ۀ��@�aCNi���P�
#\ِ���,7��P9�26:T�5�	/���\��Ss�H)����McA���Ua!ys2k�����ռ͉D�g&N
Qb3r���-bz� ����go-N;B�����D]��^g�C�4�G �>�b#����.#�z����]$m��]ak����ӟN@�8i0�.���b���uK~�(?�+@j��r:�\��t�H���Y���?Ȫ�V���H�(Җ�&zm��=�{��9�P$q�f�>���9�F�rPtx���H�FNu����)7��H�w�q.�]��m9��r�����}iVf�k�yN\�d���/Ҙ=.�|԰G�)!�h���6�M����1۰둞�.8��ߒ�t֊�if�+��X�E�91w��lP������?&p�[��y0A�4F�{�l�a@*�t*�9�L{�ˣ�	��Ocb�3��!�u/��#g/���=�[�GTV+7!EFy#�el�6�hܴ�=J囇�B�@�;�l�`��!�O>e[$�\>��Y��W��ܻ�U�����#g��mw�)9]�;��9�:�=����S�������k�T�"��o%�d �K'-頚^���	X��EB��H,:9�Z�-=v�O]��V��?�.�_Hj؆v3�1zV��tc(��?�M:�p�j�4���ԷO�[]T'�Ч����\n��Y�S�j��V:ٴ��=e
]f�����»(���*��U.�gH��8�
�@NUz�jq���E�K@��G�ј�ΡنeT�C�
���i)ɟN��&G���/~ǑH0*��r9A�d^ò�o�T��b��=��e�0�Χ'�$є�xR��E�@/���䦧��w�
!S��Ѕey�Efn�ÿ�D@��QS�� ��U��Hn��a�����	m��"x�#�dc&Gn�yN����q~�)������!���nyw{)@m �,�]�\���lAɉjM �̑��E�K�X*��c}��WX&�C���+�x�f�!iK�P{ϼVI�]E F|���w�0>���mOrG�
)�_e�x��c>����������[O����/�L�ί%D�1׼]F�t�22%�e}�)�%�1�3-���$ٱR/���F/�x����6�	���G�)���Z3^[�G�����x�|��lg�]w�6o���#w ����H%�;�Mj97%%�D��(��^��UivWX2�j�F$�W0�|�?_E���8�������q���U��B��@�SUdY��o9�i �ր\{��|��#/��U�MZ��WmgB�r1Y����I���q�}�>y�g#}n"�x���b�};9Cj'R{����ؗx+O�B6���E�L�W���6���_�}y��H4��^�x�l]A�P�܈o[��rpR�L�`����za�87�Jg��������<js��w�b#h?�oV��s�v�Z���[Q�)�����|3�� �t"�F\���=#�����{m�a��mB�]{q�J�a\c
��qg.�mF`��?����G�N�����P,H`�Lak�!V�������s�Ma.{���t��}9�T���v����`G���EV2�Ϛ	���I�`�e�ۘfړ���4!� x^L?�<]�e���)i�x�SKρ;�:�Rbv��H��d}��/�T;٣�-�t!�k�� 5��mo�����|��@8�l�wd���-4�3��)���Ng��:d���d}���F�䣆 �A��m�����_7���A�I^���L���`�#n+\�b�*'ä_ȟy�_��4A�$�]���OUK�\p,�j>�������Ċ�8�d�i^`I;��T?��s%`8�g�0�y�$B�S��S.�n�xɸ�-�[��_8@�!�Zq��}��*8֨w�q�R��z���3��Ө�.3����xf�i�!5��75֓��M�H�I.Lf�h���-�Ҵ���K�Rbf�$J��.T�r(|3&�!��f}�$�K�Fdn�_Lf��'��׸	����EC�������U�m;eZm�'�K,�9�i��H�j��p��Au����6zԪ��?Z3�ʂ�ݍ�P�f�kw"��:*I�j$�e5Zp9s�y4r��fa#����/'�|��=��P4�7&ꏩ`Uz������/*��Dа �HB*��9��3��(�<��K�a7�خ������6�/ɝ��s�6m%E�F�ۦ/����%�7l!;�{m�؎/��h���t��ޭCce<�'�[��(l�M���yXM��f�O��3ؽqKD��&9pBJ�=Y^��U�#���~%������u�� ��M���ۖ�Y�ú̺vo�w��� ���fw�T�����"����Z�	���­��o�e���~�T�gם�Zk��
�[ݲ��l��)9q��zm�p8C�I��i74P��z�J��5Uk
y\�.n{�ON�89*�M.e���
Ծ��Ơd2���D^B�n��*��p%�T���X�8���H	��9�9|�N* �o�{�N_��_`������]��@:O�4n)�'��u��NJ��ĕ�-��T7"JVU�^wōC��De�ՍT��T������b���E_���!�P"E�`��k'@nWh
@0�*�S7vt����/�a�tV�妱cqv��i��1�umY��:�0&{��}���e���J����r�NNd�8��.�EVN0r#
�����SK�R�L�^"�W�ύ�:�jl��U�������~�1z�*�i� ���@ 6[ό��@
��)f=b����|��0� ���2c��J��q<�Yc�R[y�]�;qa|��F]���2l��2�=����$�K*�d:�ά��PQ+d�H1w�x�B�LQ�;��4"�Z��L�U��Bj�4A��`�������ex["mE����	���L7LV���2�D�xC+1=�~f��ݴ}�ȋfXpG]�����@�r��7�8��M���o�_]���J�^��S��Y����7�d=.���˪���K�ۃU�l���Չ:��-�s�����YUR��r��Â���j����`;`y�.��A� �e�^<��0"�� a�"����p��z;Ʃ�!�B +�H��X�C�x^Y�l�/���r��&ص��*�u���2�*_j��Qبhve}#1t�e�k�Z7�?�KXj�բ&7)LX�$R��M��5���&2��OGxԏ��������Th�>���xF
�g�ي=���If�)'kM��O��i�3�<���l&"䦑���6J�s"�S���_P�$��D@���é�љo�`�L������K�	m���	^��o�Nq��Gֳ���He�X L�;�St?L��8a"S)2�j��ʯD�bY���{�+���$�Ӛa��Y�t�����H�f���'��f���#~�Ke���3٘����o/�r-\"	Կ��Cz���K~�bG�MoT�Z��/c�$u���1
K�?ȈF%ǤIؾf��to�ߔ-�o���U��&P�֩l��7��r����QD`�#�5a�������#da�+ӆ9A����u䚞���k��p�+���=��Kf�9�����]��Q2��S�g~)C���8Gw����߿�6L��g[=��A.MBb�jT��c�:�
_�͈�j:��.��Dk4��Zc�ߡ��w 2�f[`�	1�L��	eʀV�j2��m��<���8ҥMR�J�nm�܈��8��Ol� ��?�)>
��,-0�j�i�*dtG4�lb���8?H�����lP��]��o�j�{Q�2�ϑOV�7��f�,Dʈz挷E?�z�|�|�8� pԆ�ȩu� �UI\�T�F�Ő��@��Tl<�x�5$���q�E��V�le�C��ln�8�F�:5��𔝭�I5-��À��n.?I.��)�
ɾ9��B21������ �&��!�N�*�*� x3� �� �Qm�/����s%��WX��eoA����WcMw��Lc��317((�BW����$̆���z4�w:�Ԡ>��FÚ��dZG��1j�����5����e�B̌�_=k�+���?�v�h-�WG��z���V1��\�ׄ��>�5�ܖA��zru����W�2#��X���������ͬ_4��&��a��b��8)7y��l{�YSv~�0��ʒײ��/��,��T����0
L�j�Ӟ��p�
���IP~UJ+@�ywd,]Ub|g�KG�F
l�,:(�8Xe3Gs���`�.��K�@qMR��I�����.�g0�g�W��w�^����֐=�l��������Dិ���8@@�A�`Uf�"h���e��-_sX���"��*�z�G
���W����-B�%-	�ql�������H��H1�����p�Wd�Il���YarD4;����/��@�,%6@�9Qq��(���MD��`A�s�CY)�y�{��ŶD%�ݩ��g0��-�7�:	���	jg�G�s���4��?q�O�_�N:.�L8G)���t�&ˏ�7�5NnZ~�0�s�$`�Q���g��V5oBfP�)σ@��5_
Oe-,bբ�j������u�p:l�,�0>��f������s��2~v[����f��z�NJ��֧�L���ڜH>�J��H��U��L�N�p���t���֜3z2�ig�j|�\��0��h�W[WFp|C��5>��r2�e��p��=��o��\EC�u�Z�M M�#R�zm���ي&����e�n|��$�M�e�Zf���ȩ����h�jl1�J�X�K�JJ^T��;�7�\�(ntF! }���氼���l�o�b6���#�v��v�~�i�`!,[�V�<���&9}	��D�`�ND�h�Şsߕ4|�uh�e�x>Q�R���t�:�j#����w����<?!.��@8hr�{@��a�C�Q>�"9B���I=�t���xO��5o�v�[�8-�s�H�;�yߊ�� �����B�'��'�8�c�ޛ{����A�- �FzN���jN���� [�P� p~XC�V�I����i��^C��Xd���؅�sc���h1:��^��JD���ki>�v��[���ؖU��E���lk[�o��"-���W�R�gfK?�k��縈E�f�c^�F����CE�S޺
ҳ�����DS�fFC[�+�_�gN�kl)˳�M5��ύ`� M���)WQuQ����t�g�W��nOSύY5�;��)T���C�;�g���F�K�7�t4��0(�y�"���H0�#߭�t삏�(�~t:E�	�J��4��Kh(��| /{�w��޳)9���֯oj~<@!RE�ȍ���Xi/���O�������0P�9�!!OE��*`as���U�MX� �b��3�B8̂0Urz�J:�����(l�ȏU��s�Y��b�U�0	�����4D4:c(P�qNHd*n�|�@�M����&~���r��&�v�@���S�H�=a�%n��~��UM����̦�%W6*��I�ѣW'�ڔ����l�j�r��?��
�D;�r�~�-.	n~eh��]�(��<�U�0��r�h� LrS*��bg�D/׉��,�.[ ���r�*��>z�/���-�w�V��W��2��5�m���k
�u$�� q',B��KBM��e���5�?����|ρɨ�KV X� /V�`��K}�˪��W~�E�#;�z-'O��m�>>���lؐ-�ς ��4*�q�o��ٶ���Yޟ4��5����&����\:���DU�}�FM�qS�0�]i��2[9��|C��F�)�#Fe��x=���S��Y�Q)���sPVJ%�%^�|�����CGom��x_��"��6+���H��[I�������e���]����NZ��O�
�����ܒ9CQ����i�J1�������3V�-3�b�h}21���N�0��֢<��|
�z<���C�7�쨈B�-蝇G�8�����C��!_�]��7��2H�p4�eu�v�;ˠ
�p�x��R���	�*��x���6��<��D��~�
ū(�S��㶑���ijOmW��(#9V���5gQJ���Y ��7�ܞ�l@�)rS�r[H�ilv:Q��5��m����^��z�W�&J��At82'{:Qb/�IQ�O��z=
I<�/>�!�I�о�ѭ�H�&���H��h���=d-���mP!���I�v��(�*V�aP��H�X�mJ9�\'�6�E�U
8��5�:�n�B[M5���t�L_gXu�1!ڞq�;������pRS�-�w����s��QsK��YLXG���v��%��ע�_�!���o�F���.'[I�]��]x*�zW�Պ��IN���!��̝�l�Q�@��e<������ÚS�T��p�a��P� ����V�u�d��O����"������aQ��G?� s25�캎�[Ab�'sP5��J�.�����,	��S4�E)ꉪ��D4�d�1$�F��*w�a1��bß�߇����*�U��>{��]��R$NG@M��p�gb����Fw�ek;j-�z���;�+5-���`1].�v��h��1�6�q8�(Q�v	�Aɡ��bh����s����}l�G�;�j[��6�v�-F�H��W�N�,�1�y���uc��E�-���!�Y&c�p������R߸�Rp=��}5 q �Y���K���5�>'��5�(Me���f��y�7��O��CC%��S����[=�x��T
�${�e�PE�A��Tk��Ml��11���c����\
��1?X����)g��ؐp��h�J����K� �o�$�30�����l��D<B�mɽ�kO3ϱ�P4�p��w-ﾋ��k�(���S��#��
bўww
aT�K E��I,�C�nY�_e>�n�Ņi��~������{�ca��FRR|OϘS+����	��CD�C��n�����h�WP��^u��;ޝj��UD�d�I*D�1ݺ�j��y�:�G��d���7���zI��t�g�f5�([��3¾S5!�l��4 �&:��L+��'�_�o�N�z�Y�(����,��k嘧���H`h"��@���ClSp;���*j��ܥ%M����Z��ɕ6	��/T|]0Bp�NM�kW��X�w�������y��R�Z����0��)�T�R�9T%&U.߬�	!4#X����$G�OŪGk���k(h�M�(�jd�F��]�!h���,�g!|��z�_�Ϋ���H�nX�U���q��˰��Ԑ��v�H�Ҵ��s��Ia䒂PhI+"'>Ӳ���ƟM)tN�Dt�B,CJ.��$�z�G�y�K�Kۏ6�˝�n�8��`׻�j�#�˯~�
K�d�E��	� �ڜ?���O��< �Eἕz�PwRK�p<���Qj�0p�I��I �q5�7�����j�C�g��������)}���p젌��N�1<hD�+*������$��彀H��d��{��4�A��ֻ�p�A�[� �既5l]�I#c#i�L��8��M�5��M�.�ܤ蓌�t����q�O���t;_Gx��"\
���΅�B� �ݴ[ry�[Tb�m�<u���D�E
�3�P��l�N7��]�&��	��-����i��e�z��?��װ�
� �W��.�}�A�!Ob�`e?,d\Z�C��B��;O޾T��H�,���`;h�'C,�E��&�R�ǳr�qLͱi�Փ����������V�;+�Û��=�P���[kq���z����H�c�
2H��N ku���4r1�җcm<������χ�.��p��G�l�6��(��C����䃈�6�?	_M��|��0+e^c�C��9tIp'��o�����tA߫��sm��̬�E*]��Ʃ!��s�P��H�����#)e��B[����u�]1�Xz�^3Z��m�>���R��v:=��v�~�g�)�Q�<��˨����������xk��M/��+F$D-�� ��7�ˡ�{$}�+:�/��h�����~���y|Ra}�^�� q#JlH+� �3����4�����v*�'���J��*Pӡ3^F�W�m7��nB�}/{G�+b�2�I|9��i���蜷G��zV�')�F�.rm��̓��)�@�	��F�B�t^� %3�����ZDsJ�Ķ�����N���>��x��.������FB�����ο�z#��ԤJ�P�N�)a���K*��#���\ԽH�`�<�����6��چS�L[����5h��6oCx3	VOh�z1(�ǖ^�5�˧�Hy�2��k�%f�5����M���p؟�-q�[&E��B�4���C�<�m� [��:O\�hJ������#]H�ܓ��N8ȡ�^I�Q��i1����y ����|���y���
�ks�@��|�.C��ul��:/�u"�C*���N�l��z!@ e�7�:s�O[���p9�	��h��2pF�Em�Ol�=t���$)�.�b�KNț��,R,� ��z:,�m�����H:L�)�d	q��/������X�W�7jʂ8F���;�FE��n������g*��ݾ�}��R�0z�`*m��5�!
�j�p����:<��D��2�bg|!���/=S�c�0"(g�&Q�W��z $
�1�4��(ho#�(,a�^5�a�@�Q{Ecea��TXC���«L���<C��u���s5�9�Ѱ*��v�C�v�4O����63?$7[X��6�\�脔�,	�8�.�T̓�|Р��YSI���L��Kؕ���RD<�\˗<f���$�tY%�s�EGT�C�(t�>1��W�Jђv�B_��k	�u��Q�v��bAy��a�!�D
�*�L�ny�c�����h��د�<������%�icp~>�?Һ�po�����T�>�mn�?��6|��$?�&��q����F�αm���d
~�`�YC�0I9�M��v5�1�5�i�u�J4*P�f9����V���*�4e�B�d�}ϸZM��/�q3�3�ܙ;�x��ˣ�� ���Y@7}	X�<Ѷ�
��51���"r!�/ӽ�giP1�{�`��t�мڔ�c+�8�)�_!�v��C��;����<z��`�@1������6#;D�s� ��zg�� ��y�א�1�;���V6Jq)J�@��vbӀ"����7�)��p�F#Z�ܜA-p���:��7�+�~ll�������%�",b3�M�|��$���{7(	N>H
�Y��$iW�hJ¦:r����F74\���m�|3���(��V�/}��Y�}�,E�kۤiX?=�*�-�]��eDF��T -��e�q;H��������'� J����с�C�j�MPxi�a�3��5���_YoC"�㗬:�0�e���#����\�ܔ�ƾa����`}�6:-s���};p�<�����jݤw���{�bG[T��i���o-ތ�#�m�9�X��iad,�Q����\��2Ǧv��#�m
�@�SA���./�ֳR�kf�6U�nĊ.�<��e���I>�ٛvp��#k�����/�D�攁8册@T���_� F���-:�w���p��g�g�ڴ�'�6��ќF��-١Y����p"r�����3��C[�H���޹���ȋMg���Up��xG:G82P�4�
t��* �c�5?h��C�8�9��oq����ҕ8�	Uؖ�Wͻ�O��{t����{i����$�M����*�i��)B���m�d!��uןZ����*/L2,%��wN�VQ]Ԩ��;��!��p�g��=*V��؅9�h;���ٵO.+%�+[�a�%�cu��1ײ�%@�#��a�8z��kԏ�W����7LmL-�k)jX�Q��$���OD]A?_2sd}De���F�9����oU0`�6�氎:�����~0}����z�����o� ��q'�U�%#j��V�l:-��j�%�P�s��zy�wO!���Jc�1������E��@�QŋmPU��V!t�qvj�:��f>m��h�p�;r9��(�`�Ac5������U5����D�,H�CX�êe�LOU��J��Eu>�����pl�S�ԧNR,�2F}�׆.MC>��3@Ϊ9Ũvo������~Y?qQډk�'!~�^Dw"�R��'ާY�?'f&E�W$�.��3v]�w��j]�՚\��8��&%W殑U+�S���>(z�T��8��o�2h�}k��\~�? �np�k��MX��.��[���j�A�����=a-7��-��숴�?��W�g�Pa_��E���Q��������w��3/��Aͭ�ƥ�&��V "�]��7F�9��"=�6�\!N![bB�^��x]�|����t��gx'3(�l���.�=�̚f�4����,R��8�GV�#��K.]���TD�.U� zY	rh��9�h�u��_PW=�_q
��o����ӘEQ��j	z��w\eL�����jyy��w}�W�8�S�=ţR�g�l��S�G��
K]��������<(�R@T?��#f�H��3���gq�\Fbґ<�s7���˞��+��?�Z���>��:��n�����cH�����"���&�D��8�����f�)=�e�{���q&����Ÿ���"�v)��b ^NL�����>!�8�GY�g�$�Uڤ�W��!׷�`��Ȉ���C�e�K�#kP�Z��!�����?��'��LE$�b�N_���L3d�'Z
�ޙ2��!�eO?'�U�����1�(�tT�lS�O�8��}�R��j���v� �ӑ�.�%:�qY Y��8=�X��H�W,��=��,ߌj���w������:����H)n�
�֏�?�JgB.���E�`w������՚�7�����᪔� �6q,�&�54��h���4#�^�Ю�,z�1�4��Jy��9��L�0�r�ए0k�.�p�v�\��eJ��?�2�8Zc����	����R��Fk8�p����ؒ3����,pd�@�y�:�ڻ�r��蘜�l�X	O����1M�eA�����e�걍��t�s�~�#̾��@@B�*��5�)ǔ�4�hͅE�\�Z�{o��a&!yA+��^�/ZSɥ����;T0�u�q�)�	9��	����^"^�?;��a�J��,=4Ï����y14�$��|��;$me056gJ�q?Ӭ���O�G��5)L�lj��۾�CW�?�O��]�������_{g��֘1�$Nʛ�<�GEv���;��;R�uP)+��zU���7%`k4kk;��r6�u`�;Rq\C�g7AW�=�z,[�a��왌1�A� ��g��}����]ub�4�3��pi�ŕ���3d���%3j?{#4�E��EDjz�c�s�7L�}��9:���sA��.Yױ�h|�;m���l>0		q<��wi+x ��W�ջ��ɬ2��a�ʅ�Ǽ*`u�J�M�a�I��;��d~�g߈���pnE^��c_ډ�P��bP�]��FN"Ѽ�յ�(����T��Yt-�$�U�o8��s!�CU�O�,˘��8gi�����8���ĥ_g�o��d�H4�.����\3V�0�B7F- p(HC��4���z�ͫ���݉|Yک��̊s��K��?��I�Y�`O��-�|dGe��^vB��n�ls���_Pc�v$19�Oٯ!~�8�S��Ӌ��*Q3M<VR�c����/���f�:~'w?��ُg�|��#l֒�� �;�OCdH@F���h�6�d+Ȧ6}z���l�I�9�	~��m�º{W\�#]~��wU�DG��΁����j1�x�
J��LsnpK/B�A�/�S�-T��V�f�>��*�?3�v;�L����� ݙ��C[�T.�B�wm�"�埣Mu�a�+���0��"�i��o���8�����4@[���jm_S����OhC��^n�K��Y?aFy'�rڬ��<������Z��&�F���rs��Td�\3�����U͐s�'��ڢ"���¤�-s�k��6��6�rs�������W;D�X{�,��
�'��!?پ8�|B65�dYY�E����D���ʲ���l�F`c�o����h�2����bBH���������UH�QL���g�;9�j�i���i8�L?�_�ç?��@a���#���Q�J#���yKWm	Ԥ����_��1�����zI ����n��!&y ��G�Mq��wW����� �ښ�|z{�pB��dw��a(�%�5�Laf\��d�$4U�(��xx������E�p�RO�*�`��X|�>	3�v�5\���z[A�5�b�rDv�8�]�zCіtc�{O�B,�1h�& ��F�:^T;��MB1�Z?�؞���wᙟ������^okJ,��wܕ�d!=/n��"B�V���N�辎3���4	��\�x����W_��+�dL�j�R^umz�˛{��Α�`��R(���`���.���l��.V��jǎi�;/�sw�����X��`��%,��_�y�ܯc���v~f܁�(b&R0OE�G�'"��"�~�6"�r���o�w�Y���r��M�qŗW��B ��� T/Ja�J���:�Q�P�*>҅GK���)���5�e���Z:Y�.ziv.��DV�6����o��]�51q=ݻ��J[FJ�X����"����{��3W�.��m�mh�iɸd��h.������|�mS~�M��ݸY�jҙ#�A��0�g4�ޮ�^|E����N�Um�k#Ԧ�6��:f�0Ξ����9K}?�a�P��Zv�ׯ�-�2�Ϭ-��D�`4=���t-S!������7�`�(/��l�,�6�,ւ�;.m�I�����[�am\�����/��l!���I&��b��c�0�W�$c�W�h�! \������H�`!ǒ�������0|���L&޲�V�/��?>�I�w�^�-���&e	�?�$N��|Ԡ?It��<D}%�5�l�}�}�"��XE��g����E�6A��(��6��E5���"��/���ca���;Y�~�Mt?�x%ɯ��\@�aq,*b3��]��p��mF��yT��V�ݣ��1R�����Q���Φ��ǻNn �n��d��wܳĘ�Q�bvW:[�1��渖�W���aڵ���Ѳm�d�r�#�g�݊���t�:5�]��Q�ݟ/T����)W�����>y�5��B����pke=�:�Bt���W�����O�W��S��b��K�5s�Y�*x��Jh�Γ��^%XL�urcn��&GW?s�=џyz�	l�n�w/�	��xz�vn���AD>�%�i�$�P@���PƩʺ��;V�7/̵���w��I=�tE�Ne-����K��$	~g��S4���N�'ѝų�k!�8 �Fh����ع!��H�^���)�Q�:���"��#�W�VL�T~X��bX
;_#EMF�&B[��(E�����ӪF�N(��|LHN�u��Rߋ��{@�m���D�HY�X���I\�S�W^��ê,�ٷ�3q	� ޟ�-z˓�tٮF�]: �1�:g��O����+}�� 3��W#6�ںD�������o)T���Z�d��q!��P�.���f����5X��?\#9ϣ=G�!7~
��ҽ"'S�r�����k��!}^�=�*��f<ԢE2I1�x�G��ƪIn���=�LC�!����f2a+۽�zT^�=D�����ِ�ᨫ.��aØG%]��0����·�َU����ba�7���<p9	��<JG'��ۓ�b;O*�ҿ~hgH]�A�{�k?�j��
�p�К��;X{1�=���n#sU�2�tZDF0�R�{k��h�ExF!���?�����;�s�/���oJ��5N���6�V� Gt�t�u���?�J|��ו�����&#{46�cܜ����ĺ����*��O��`��l9?��s��]���HA7����i�y�E���}�)!��-����sH(�lTrbݿ�h'��Aqh��V�v�#���}96{5�;�X�m�4���RJ������1wa��2��>��"ˁRk��HH�S���{����&x�u��؀�0�쨨m��f����hE� KƋ�J��@�?$��.�v�iU��>q}�q�L$`FV,��F���: [*���Z�i�MAc�Q����)��ND�W��H����ʌMq������-q1����P����,��EZ�Q�R��DD�/s.��9
~�L%TyCoV��}�.�VTˮ���.ۅ����6/�[�맀�$���C1���@�j������|���Ӡ��::%��k�9���Z�O���/é'X�M]^e�{v�O<?I$�S��
a�1(�%O���ݿߕҿj=e���M�p�<���g�}�c��-B����AIj~jD�s�D-ْ.�yav�k��q!�5	��������}�Z�q�ڋH�O�����W�5 H�5�<,ՙ�\���Ղ��f���H�d���{<V��Z.^�4��Oρ=MXi�\�AʌC����������jZ���w�/��S�{� ��X�b��1�.
��2P������g��p9����^U���V�搑�i��c�ۚ�u���AlǼ�l�aT� ����ĴI��I�;� �Px�h�BQ��\0jeϭ�³�wG,[�rU��~#��7-��w>Ż-8S$���8X�%��	�M3TCvy�۷�Zl�K{q[��U|��>]��nt$U���dU�k�#3�vB��t��_k�����B`�o���	n�+hK-9���bbv���CO���S�	C�XC�s����x<��B�Q�����:񤠵넕>�>8:�����2S*� �H�`����vnx�\���&״8���Bkr��sB,q�	"�i:�����샂�6L�Д��γt�$œh�SL��������������kڕ�͊OчA?���I-��[)!�55n�q�F�ǃ�4��@z T�'�����ۗP�����늞+�߷R?�	�+p^�O�"���>��T�6��ٮ��~V�b!�� z,$�1z�;�bC7��Z̢
� W��@��
Q��Ks6�\up��F�k��o�1����[�c� aw��`�?����3��
_c��z�V_ԆPY+	_�ҩ�ێR���|���~5���c)�����^�~GR�?����J�Ł�r$C_�"�6ќI�>��4<80��1����/+[ �M	_�y7FYS��S�I `��ݬ��4����t� �| ��I�C���/
/�z,�}H���%�8]h����������R�]�����G�{�4��]?�f`��nf������q<�<����hv��^9z����C��4:�NEƄ���z��t�C�蝫�qpW�-mֱe��d�T�We�P�kf#�9�'�'�2֡���Y�%�
lO�'��L*�Z�ZuN������uɮ8щ)C)����ʔ�>i�X_�o�I"ck೘&x	�|B9`O
��S���Q"�\mK��ŦS��q�8�1j
�x�J��4KYU��eC�����7�x
k�aVZF�;#�+6�會j�J+{o��ƽ�������ط�u�wj�Q`�fԿܗ�>�%52��6{�����苅ⲜNeU#�FNnŊW���,
K�B��>Ϛ%H��)=���l_�qM�-h��[�*��=��mŰѠ�6X�ȩo4K����E;�����p��l���R�?�uL���k���@����Xo��z�k%��We�P���ryt��E��]�A�M����グ�X�>��	I�Y��L�X�!��FFtS���A$�;&V8Ic*ۧ��-��`�U�yW@j씸֤P-!L9-�#�*��ǃ���Gc2�:��^�=�3�U���,����Q~x�X�a�}���(N���80���%^���
|M��u���wbs�먼��1 ���V��"HǛ�1N� G#��������Zxx3HSC9��<���ʒ_����b�~��Q�#p	���#�ma�%ܲT��p{9��m�J�_yD��WC�����E>z'���ɜ�m-5�sq�)|�ߕ(�Fȁ���0����d�������󴥓�Zh�a*�?Fs�M(_"�Q��	H![���(5���3���,�Z����)�����t�Z�1[܅�Ԍ��ľ$Q�����R��D`�P��?��M�|L���w�s�#˂����@:���H����l4Z]� !�K�ጘ5��V����փ�7�t[��j�`�
3��a��~3QC�ot���;��+Ҭ r>��P��N�^m���(������W��K[�:�h�
CtT�9�켠�-�]�5+$���ȍ=��WCV.?�i6t����N�sz33���
ڛs�a��*�gX0��'�ȗ��r��'��S|%�*��@j����_Y��v�S��E
4�N�i����.u!sG�*�'�����Dw��K����e���~��Lm�k�z���&y���tww�NgP��j������HeZ�yc�l��'nz~X�)$�݄ *=�پ�KQ
�L�Յ���Χo(C�p���9���o�I��)E�;��%@?�U�A
�{���x�=s�k A_�}c����3
Kn�:����򠔲��1Kh�����ZF�P��s���1���#�����P����Ԭ@6�6�l<� M�#���dϵ%2�qh���ЭVab��&����x�=eS�zmҨ7d��4ll'Z���Xw��?�N�{�&��T2�
�Q��i6�$���o�k�q!�ѕ��r�Pj����x��[�&��b�'�ʡ���v�E\�j!���Z���&��ց�����D�� (*��?�=��Dh�fpDo�`�/����iٌ��5}0��L}bM/�m`�T��,m�/�O' wp�����������m�P*P!���n�����x`��=f�=����S�ﲂ�E���(�6�*k�B��'BU?�Ld�O�Q��
m�.�~�S|��o7��[���:��mX6��׉o07~�� H��O�WsX;��4�)nH��V����;�1�AN��,Jա�F��U����������H5�N��USN�Hb�k����`�QC�o/�]v����1�IZd("rV�H��u}�/��O�ձh���}z�!}`1�W���Q�AA�Eb0z��8�rM0߸�$�v�PW��Q\�8�l�v�Z�M�?)����.}��r_����b ΤUJo�^:���H�kI߃�%�҉,zz�=a)-��]��O�����%��̇���A(S�F@I�h����ކ#4��W@�p.7Y#�S�D#�K��,�k0"�c�E�e{�M�"��5ݼ���h#@����Y ���?��V#%����"�s�)�"�7r�E|d��H��� �%�F�v)�;���QRE�b!^CV�.�|ILgM�<07ADt6���IK,�~v*�ک+�5���h ��񖦆;m`���$��	d����M7����e���q��[r�Cé���L�f|��,[Kb��NiK;�Y^�^�%�2Ӂ�8�s.`��H�$jf�̄���>%�E�a_�G�-oQa�y/ �)�ԣ���N$+��h�I �bL�Ml�8$-@�?�>��
��>���\X^0`q�IKH� �Nߚ'�*�0R��M.ȷa��x�`R���v���	�5%�M��*c!�����hq
J�Y�|��TA��':\H�e6��a�N�W�|����p�a�i!)l��V	��{��WV-᤮4=�e�_��^�@.���x��9�@�\=���t�K�����{�h_$]�]H ����K�^���TC��( �ɵ��%h�Fv��w�MD�{��6�p&N�rg�~��'�'��u�]o�ǉ\;ZU�լD�qO6��1���;i��i֥rZ �D���?O�$Z�L=������l��W���-��_BE��p��	�@��֋m*��P��k��Z��v��"M�t�Tg}F�Gݤʲ+��:*%y$�"��n춁z���i��h�!���v�C͡����q���ۧ���mڈ�=�Ϫ/ *��)�ѓ^������ [�VVs�����]�l�q�#���[�F��0�^l�oO�z���x3˚�B��$���E�oś? �e������LĮ 7;X����Y�Y�X$̺�Lz��r˂�!t��Y�քf�o��QB�0�H�^�+����|���	T�A����6�/�(�x���#�#6ܣWdj�7Q޲e<��*��T@���t�QE2Un��{�[�̌".�8��&�2PH3!�~�Ͼ�/���L��E8��b��O�ϣ�ep���q3T�?hh��>rچ��Ip�h�#�i���"4ܦ^��ǜ�,��a���W�i���k��t6��B�=��HKfU���tw���8��hg[�/��*?8�=_�!������'_�toK�� �7��C�vgL���?�*N��S� ��J�O�ZR� 	��V�$��~���&�v�U�w2�}����h��V� P�-�Jz�� `W�Y����4*�"eN����?����N���u�]���$�u� �0q�K��4�f%�������s`�L��;X:ww��6��o6G���ߐ����s	F:�:������K����K㏘=vw��j�\��74�$J��� =9ђ*;�VX�����p/�'k柈�U���BQ���#���L*�Z����t���0��X��4[*��Uj	��\�m����]��vz�����0���z� ��(���ֹٰ ��7difi�fy�K�3^�B<�t󥪨���b�ljl�r�t�R����.�����N����cָ��n�!
C�W@e�TV�ٚS����3�����:_� b=CS�A�~�X���=���/�3��~ g�Ҫ�bUZw�-a���契���di�o��x���/�%gB�c�J����ˈ(���D���,���?&io`Ǿ�l����5�5�?�������\7�L%&��J�&8�u!X\�-��IX,�wen�x�/�G�E*+s��(�^�o����_�I����Y"M�]�{Ynw���t�Yٲ�b��-��q��jC�"�%�Z��/x�s�Y����	��OP^!�~�ǉo�j8�b���?�c=�n�h{k�&����]��n���N@<y5��b��X�u�[IP	*E�j������-^�LP ��t������G�Qjl��xR��r��1ѺV�PГ�=�����m�t�L��(���r >�bT�!��wU
�)��~H[6��&n�jڊ�a�/%E�`��	j�Z.1�C�L���|^�XXTx���8�
�7(st�V���v0���y;��E#
j�
����	!�o�|;��X>��͠�G=�A�X27�J��k[i	�M��!�WI��1(�����0�� !�qv�f�q��ۥe�x�ڼ�F�̠�l����t�2�'X���qh@!x9Wp�yı�Sq:Ç��
�Vǖ��J*Gɯ�f�xc(���W|�������Q��fo���F-͏������Z��J�z���m�C*P���4w�hS�����<�e���r�׉������5���0	���h�&����!�|s�H}X��
C,�w��&0�b�?��~��=Vd���^K�}W���=��:��3@�[#Z�)n�?�H���s�8�.� Z�cS!�|j�oÓ�xh_�
>����c�"4�ĂDu�����,���3�GYY$� {-�Y!�sx��@T�<���$���J���ԩ��u���<ހ��/�G����?�*�#�(6��_�?Z�����M���̵.;(��G�d25�}6TZ˼Y�4��Yf-��c#UH����ɔ����2p��{���a�a�n��@�H�Bp���x��o�ǈfYs����8��k?��rN����ܿxRu�v���w�wYZ!u?kַ�ɮ9e��m�7��t�����#%-�׃}��R��5�K�k�F�!%ζ2Sȱ�)�$��ʨh8ڰ�-�D "�ض3&�;�x��X��)LQ]¥����35�6��i��B�ѷVy�v�i��C��9B2
a�ߎ$�|)f�,�k\���t��=��6,Hz���ĭB�qZՋ:��c�Tc>�%m(@ۈa�-v������ђ?wjPJ���AJP�<	�q�����L�r
ϜYj���Wj�w?յ]��5%�B�ܘs��`��:�x���e��!�������6y�|b�)����ێD�m��YW]Ds�s����N V��A0���Z�_#��ÖV�zs�4>�����֎}��ۂ$���JC��2���m��^�_�f� ��%�ۨ�D㯩�Y���Ե��0EwxY�9���]c�5�d�V«8t~ԇ?��h�p��:�`��i�����ǝ��KU=/M?��&���*Pв�0�����ރ����OW���;�Y�XCVߓN��U�#g�E�v��"�	hQ�� �l�9n�FS0���yh��.0˙�G�і�l,��>�ٟ����N�0�^8��5ˇ�DacV�e��Q��Z�e�ɠ){
B{�U JF�HP/��0/ �}:$N�� |x:��%���F�Qs���lV��W�����3�����Mq�͆����hL;�5gn�3��=�&��b
`��5�h1B�7���#�or1��?Q��򽞩󽛐�H�y�`;�E=�Z�C1��H f;c�Wot�l!�KQ�y��VO�\$�`>�Fܻ�
�%P7!l9�����dT��˔���/f���0�^��9�O"c��#�q{�u'�a���8�/ !�mc�W�G�l<����3oQwS}B�I�� f�9�:�aI7�i?��w逮f5}��f�V�z�_�[칥��g�PM��y��!ݭBr ���)�x޾�ǵF��jVT�h4�1hԅ}�-G���f�)�<�2�)r��Ą#2M���M��{n�����x����gU����)�#[�6}'�>Px�|o������%�N>U/|q�-z��@&WP*G���2�m�F<R��O�&�U�4�oUƱ�EK�/KO��-��
���Ѐ�.m��ZM�!�6�V�A��c�m�����g;�4�)��b����,cd7-��G��bƓ���^�R������юզ��b���\�����d}FP�+jJ��6�@­���x�| @|V�(��N-���_���#��h�dKyRڡ'��~�oM2��yl��	�6J��Ȓ���n���@6ou�E�V��o� >�v2�3(]mS閖�9����|�#�;�g���˨Q����	iѴ��'�D%��OK�U�d( �q�w��!t�n����S�)Z�Չ���%{yˬF^n�ړn� Zk�}��7F.����5�T��K������Q��G}FE����>�χA$N.�6����m�@��`�Ñ�[�It��J�H�����2Зg�F)��`L�v*�J!mͯc!ϧzC�O;Oǫ�2�:�{sԱ��EQ�iwn��@�����do���M�KH���[����^�p�����Q_�Qڦ �Lj��W	�B���Vg._����%gAj�|�'�5q�<?�{�b����u%B��	=�'F���眧vA�=\�����;T��6��L4uP��
�~��� �&_��j���I��i�K	Je���|n�vc�S����@%?H���"g�,?�8)�m ��@����G�ә�8��:�d�>�Um�������o���Xi�v����+z���d��D>��t�K��	��ꑦ�;�� ��c�-����a��U�ء�,� \t��� w;m��(�[z�08#y<��s����]�	ʗ>�m�P�x>6�?��1�1�,�  IW\f��W���xBx���Q<'=�^����h��[��3у�~Ch�Dy��}e���c�ʰj#�G^X���沷lP��x�y~g�n�����ո6��e0�5@G�F#�κ槺<y	w&�/��{�p�� �P�y¥g9��g���Hu8�*aڢ[՟A���?Iq��3�,5�g�Φ�m�+��ې��Q�%-CqN�3���KE���n�b�Iz�^����c��;���D$v��$=���a�%��f+T�+�.+���Fn��NQ	�=�da�G<��d�1�H����e!Z�C�vi���O~�N���o_W��+�1����ݲ처�ym�����\�swY���h�^U�o��	�"p���A|�=�n��9�n-Q�e�,�aUc�j��i6�0o���Rw-����Kn�
���t[j)C%iqp�}G{��X�}iNxF��{� 84�"c?d� ��O���O�*�)���<1�ܙE	P�B��V�}��ʽm���C�!�ǒ9�׼uq�l���Ӫ]�\- !���i�Hs'�(;�rd����֋	�� ���������a��O��M[ˢ�M���Ji�Ɉ�Z�Z��j��\�>���1�{"�e(!�@)UԚ�+��3/W�(�݉pX=�H�B�K��7mm��QTU�8/G��ڕ���`�V����T�U��� 7�v����;�b�v_���U�*?G���/+8�1-��H.'뤷��T`��I{��W�@)�H���3:�\(v��Mk��v\k˯��2�E����Yظ���.���N�o���X�x,��f!+��΂}<~%[���2訿bU��ZB�jy�+�HGh�w�C�p��ٓ�?�_�l ��f���p[�<�k���7��7 �y3`T�L|RM�.f�`��b2O�����=�a��~�A��_�2�z_��+T�)����*�05��4�
�����j6�;Ey0��pUe�^� �I�	���fq�A?���1`&?�4�Ø��� �\����Y"���D]�����n��P� ������W�@H� �h�G��'�F�Ʒ�^�kx{��-ӌ�P��ǜ�o��u��'B��=�y;�J��;!u1���MOG>j6鸗*��2����K����L��X���-Bʝ'n�tՐZ�eQ���@{yM��j��k�,x�)��5��s@�q��˿��q����4�F~F@������x�"������� ZjR�e�� ֝yA�`�d��%ϓ���� �zz#	��=��\aLl�hk��'�J��O%��u��B"���澹�ˍ]��VID�i�$��F\mʠ�k崴Ή��{���e;�+�����R����rO���������MD�4 �x�w�3i��l,�C�Ƭ�3y0V�l�5W?���.2������%��N���s���]iO�U�9�Jw�����yM��H+L;w���F�Z�^4k�M8<�Ą�R73���'x�v����ŕ1�H�P��O����l�s$b�f�cG�[C�{��qPV�Xd>(@��C?�d��5i�a���Z�σJ���A`���۸����J9��qT��ׅ�{h1�(��t�mT()|��P-��ถ}���O*�ȯPi��T(M'"f��<�'93����#��5X3!�D�.�FmՀ
���{��yu=yEng��G��VO�]��y�U�U�w��*γ!L����O_R���� V�>���ɋ۱:�03�u:rc"N��D5����#��{m��.5������ـ�k�[<�xħ���͎���S�A)��'Ĩ��鬷9�->�$]g,㢙j]
 ���U�0�Hg,�X|����QpX��~�����B����#V��R9T�/�������9��	K��$.Vnt�o'����^���ֶ?�1��<ea#Ҝ�ez��{w9Ҳ��"L��9?Zsf���;�3�����t�S;�Wy>�Ai���ɍS�Z_B0��=Í�ˁI���}ܙI9����a�Ni��>'|���x���fQ�^��"ۜ����j0*P�᚝�l���g�sH8M���n��a�ܼ�-O����\@���W���`��@P��:i�����/����9�$��zBf�$;�+�tr8e�?˝�˳o}�(����|�_4���<��Q��~
�T���c��*��ޡx�����aHx�<6�5��N�x�r�	G�Z����K��S*K�ݦ<�����/�a��Y�jpk7aKY!ʺ}�ߢ��$h�h�FFH1�ݠK�ui��N��(gDg$��wP���Atܠd�U|c���_�g]Z���B�q�
���ŕ/C!{����9ӱj7DN%�rj�شF4q�dd�~-)wן�@������Ey����|�\7CeO��1fA�ݖ>��%�y�zu�t�s�=���!n��R����<N�5�^op\R�8T,vAl	��+h���ǆc�c(/��kk����u�R����Q���^c��r��{�	$�i��~3��(���V�̈l�z.s@�0x5��__b4����$q9)ߩ�A<"����,'C���}6�5~���N�6����j�[�ܠҐmEw��ݹ��	�4F�͆���JC���O�V��t�d=��蠎5�21C�IBcLb���KZy����)�{A�q[�8.�G����Z���+�x���G3�����_� ��=Ǟqz�D	��=@�b{t���u"-���z0���� �؈c'�V�#R�U'� ��B04�݄X)�8��0������fl�u�$��֕�0��Ҷ����ɹ˴�!�&g�I홬����/3�^�ke{4)���DJ�A����f%,T�!ڗ��T3f��m�GXb��ق�c2�ot�#�������D���~�� �?����c=��&�L<@�|%ܞqG����ޟ��:#/%�P��@��V�l��i2�q/�U�������U ������Y7�\�6����m�$�t㦄�Ǯ�$��$�lv�}�%�ދ�!��Xѥ���j/AӤ�E�|�o2J8E��Rǎ�P �1��?e�i���$� ܕg��w:'�[`�QY�W��/�+j~�T���nFh2T���'Y�:!G��}ʯ�d�}H���u^�
�{^�>�o`ֿ�9���x��q�g�-X]-|Bm�ף60���=�{�u7�IQ_O��ln�ķ�p[��[G��Ƅ�0V�nia�ݽ3	�������C2W��f�y�5˲�ع������a���GKQ#6 ځ��w���HH6b\�Z��;�V�V��0`�M�;UK|,��1D7J{�˿�>�-H){h)�G����K�[�>���F������IJg��	P��%���Q�{�c���AR-��	�3/�h�V��b���Te�ڴ�G�y)�7�lN�7�%{�h�9ȇ����p�
���K�5q"KIG�^�u���熍���Aۢ2�9X��K\���
&luM�:fE��4ￎ]OӬ�!������\� x����&P���j�S��T�)]�h�:.��;Ӣ�ge(jH+�|��;��経�x�O����=�����|�_�[lI�+d��:���S�. ��O�/i(�����M��X�h�sbgM�0�X�Ŭ(���Y�AE;-����yN����~�[�I�6Tn�(.���߾�3"��])���	t��?��@��,�M���'؞4Cs��s�J�(��#zf��O���H8�ś~��ٺ����ֹ�	6�xxڬ�h��t���W�0d�/
a�|>nd����*F�������{(ݲ�|��j��B�"S|�uv�k��F&u3ZY9���y�A��z���h�������C���I��?��J;Mi�v���k��?M~��)�1�Ja���91"E���4��Ս��w��S��霡)(�'m�Ó�?eZ ��!)1�_��C��@��Xp�ʒR;w�Ix./�!���/�[���f�V��ϕ��?S�G쁶�6���\w���N�i4	�kO�"��7���By,{����<���u�;�|<p�n�t����-�e傯���q�n\�"�
�N3�Sj��!�_<�E�Chj-�2֎�:s�>mu�h{�$�{�t�po���V��TNw9Cj�l�~����˥��VK�7y+�Y�ϛ�A��r,���� F�;i�1 ��˯�]�㝒��r.$ƌ����
���v��a�ɾ��G��I�@��s��m.:�	!�����@�X���4bA]��1�M8����e<n�č*ή�Oҧ���#�g���01	��������BH��٭�x�6~9��`���A��nT�򪐞�05�r� q��%z�K�(��<tC�#���&
A�ߔ¤.�m�ۇ��}!�9�ػ%7ϒ%u�<�=�o0�h�@G<4صq@���*�4����W�&	yՈ�A�}4T�<�O��$ƭ���ţY�(����@�e�f0.�ݚ�s���cO3O,պ�m*О�W�V���R�0|3g}TtϢ|5˸�{s&�H�SE�����@�o���S�����:&�/mky���jW���x"Z/�) �M|��@i�o�W�9qdK���0#��mb����$���Q���W0�M}0�X��T��.�1h��TWE�N���:��G?��亀8nMP�}�2��K+x�k�9��^p(~`\p�Q#]�)��U'��<�6ޒ�su����C�{��shG�u��S]t�t�W��?�Ϙ������׼\��)yn�em��(~�x���7�h��M#��̒��
�K����H��G�ǳ�95�Gx�e�D�\�7N�������W*�:_2˅N�n)�P�7���%ɓ�t�����<��*Fb�`�>O&�#O�<�GxB,]�b�>�����sk���^���FAN�`�S10.��L�R�Ѯ;�D�?���b̋�Q��}Jd(e�N���<�]����,�Ю1P0#��E��դA�F�+�J`�-U@�A븦�{J��c.g��T�$jR�;$w7}���|$U_��<X"�`Plc�o�b�iz�c��/�:���د8c�V�F�4co$�3�W���v�{���K��-��o��,��]� 	W�l)�iCvjȉ�V�u���T1�a?��X�ne���lAudN�uHJ��hҩ.�ě�F/�s��uIѷ�y�-ֿ�f�H���FW6/�B㚙�'{���ֺ�B�YQk��"���pDP.�T�'&;��(��@"�,{Q�6�E���7����^Ȱ��uRR��:-��^��ʕ_|�c�	*a����)R��S�������Ǵh.�V�e9�=C臰9c�ی����aZ�PLk�]y��@I�`��5�@\��s"�K���+ΰh�i���v��dL�0j��gO�߯�3�����	/5�@�'vQ�L���5�F)9]$x����ʳv!`�������)ǭ�����z��	7�~�:��y!��?��Ʒ�� }.t (���,]�(OG������Bj~��%10�Hr��m�KM�����u�$7���ۭ��i�|L�#ϣyr��Z��3��w��oF�O5VǸ��f/�M]E��4���g���m�>#��'����%����9����l�����[igt�ޜ�{v�KR������pǷ�Q�#�Өc�|�4>�N�y$���PY�����]^��{?K�zMS\�\W�$R� 6t�vY�Q�u;�|M��.V��g6"z�9�����j�����^�#�9|��2X�,^��؄xd��ݩ���&?)i�����%a���`�f�h��A1Z�Ƈ�t]q�_l�|.v���4�ʨcA!/�n����è]˨U��38�}�Ο�? �w���e�{	t/�&��y����!vE����A�N��T �O�Ǯ������X���mIV>xM|6M0\j�x?p�Y/�A"8A"��ט�4l����J���N��^�&�ʺ�O��+�n&�1K=�2�U��ӓ���O�?)0$��B��ps-a5�$$r
���-���
��K����
�RxI}<�*��H5�H�cE��m8����7}�y6�����։��h�)L�0F�ț1
b���;�j�\|Ř�UI�)���'��;��U^fg�����Jb�E���)�=��`���cs~��;a�|�J��.��樵9	�l��\ ��pWiL��֐&�$q�C8�;�^7F�OՏ�a�^o��S���BgFe:~�ʝ�����y+؂�hi����"�o��;��f~���^���&�ن͍>��-/�gVQv���iF�(,{��V��m7�~����=�۽>Nn&���B��2�"����I��VJ-`�Yƍp���Ε|(��J�<W'n;4����|"�;L8r g�� (#��
7^�o��f���j[�|�U{��� �2�֐O�K�dY#|6*�H�n@}��&�_��%>�~K~�m����k�=d	��H܈�YUA��j�!�N�\����ۗ���E,���u�
�C\1\��㩨���o�b���6Q�ȯ@L_��LY����5z��bS7T�6Y���/��p��5���-³�2�B�\?���T7�a8�&%�	�� ���x�^Ҷe[݅�G�L����?4��.�����yLC��D�wz�X�9g!�¼Yu��^9�� <@�ߑb��W�C��;��ෝ��38�M ��X�gZ���&L�6���j�1�{��{��
(.箘�bf�Y}p ��+Û+�n��m��jv1�;�"�F�&�]�x��[Kya�*>p$�j���7��2�Z
U���r��)Y�����D+�`���9X2��1N��+rk6�Dh(�kq�"�Q�+Q[R�-�1���I������_Eͮ�A��Bx2��<��\���Jd2^ߛ%�F|��\g��_��_�%����RbMS0O0����qHr�E�����2����_��H�gBB��UE@��ՇR*N0؂D���3[�R�9*�5�l�E(��	����x�p ��1[�t�_�(X-��O5�T�y�
��8h��e����~9���-s}��˴U�!}��xQ�.�v?K���FJ�T��h�~`��̷����^34wG+L������{L(ɮ6�~��y�S���:-���_N��d?�.�⠱*�\�:'���T�g�y��VX눠�ʿ^�䎀�I�d��j\���ܔm�7Կ�u̠��C 5���S��េ�S*���P���� �AP�Rm�8<!{���bc(�J�ٮ��_��+��/d{@q�����K��S!�.�.r�(��d�LXLr"�0N3�to���񼳅��u���!aۜ[�{�5J>u�P	��TZ]s���Kj�ʣ7x�uDt�9 N�߮��9u�����ԛ(�b���2Z�����Ur�M#�R]W��!��,I�M��@�#�j��Sp���������9O��@�2)�x����~9ZU�9�il4
�Uk�G3�V�Ѐ �*)�ħ����;��'�������n?�u�<B��7+� ���b��Zq��$�>�M(�CQ��x������^	��"���5��{�D��e�>^��1E |���}&�v��>�+��+�8Õ������@ʺL�\��2����Ӭ>(A����]��9Oj�`�v�Si�aS���� ����x.�q��$'<DG������ٵ��]�`*�g2�5ȼ��D4; |��|�ǳKK.�1���m�
��w�׻���!,R_*��mJZ�vʡ�gj�5������8��8J���6�k��219 ��G{�%A:�8���L2P�ɢ�@�m��/��sD���K�E��5�vBQ��2��&��k��(��8	n��Ė]lZ~Չ���xI��n���T��y~a$6��x�kM�4��H�s��ل �@�G�q��ȃbW,T-U�E0�����K�җLr q����F����G�7<\�쯄��m��E��O���u�����,���#�t>7 J���2{�Y�l?�@���m�I|j8�
�%�g�=߆���s��Q��;���EI�2-+�,~?�:��|G]$UQ�KyE~*Q��N�?���@,�+x�I�V(2�������ZJC��Sv̸`�@�h@�*�?���+��<R�����jq5=��g��fࠥ&�.�fA�$�t�T���{���t��"��
��q�R\*NkѴ�'o�y�t���wm	"?2(C������Z�o�s�A��!-ގ�	�lL
��gp{�'�/f��xhgPV�9�7���/��"���vy�>�X�i%8��{n`Qh�tNt��'1Qޠ� �����
A"hp�x:nA��+L҇�k��������"5GT�?=cMT/�qН-C�F)*7��Cg�vz���^��_m��.���Ė�W���5(��	����G�v2;��J�^
�j557\�����x�yo<X/l?��Bd+�j\ۙ�E�����1���q��hի�C��N��ɑ�����M9c���Y�γ� �_��5h)'&����d,���ф����J��m��{x���.���F5����X	�<u�����F��
� �q8"g68oX��Q���rⲅ�X�h237#0$�%f��8��k3�w:�^���ޞ��UJey���T��B<Nn��C>�3<c���(��l�
LV],Z���+t>�a�v3�M��k���D:D9>�*[џk3�V*���t1�Q��~Z�����ҫ�,ŒX���mۖ{�N"��)~�D�p?1<�3�9P�z�ENAJ&�4�V�5�hI�2�*���gU�=��I�S*/l��M����sdzϔp���B�1{�aw��C�GZɫ��?Y������(���#8�y���^��|&N���b]k���e�"��\v�*�X	��(O�&=F�rC�=��(�{7\�����n�~KJy�[�~o��&t��\�m0�Uv�_R���O&S�����u��VxDz'��Zl�0_E@���S���BbW�6K�q���(�r�����m{;�V�hd��tĔ*��?ZJh|�Pyu�!����_E���}��V�j�i����B��.������bN�L��Q�P%2�q�p�A匕�v������Oʦɭ5q�w�|��	�*"�/J{�9wY��d���p�|Q;�u�NdWpp���V��}��:����m��1��D�'Q�g7z���3�}�SO q�q����gCs0&�d+v��J;��qn�$��^n`tITO�Sy�^�`686t�@�u�E*�[�]�!@J��!DY�!�2?�z�g	R`�7��t�_l��啍�E�&Y\ �hln|�FoL���Z�A͈ �E���Z�e���N���3c|����/��mC��%l@����`;���l�N��m�B�����v&��0f"p�󈉦̓������i˱��kl�NȊ��b]H��tp,y�uG�}ۋ�l���e4��6��1�ԙ���(�������2R!����"�nvK����r*V�z @����)E޳��y�l5/$I`��S �ʧX[s�:���]�2y��h����`�k��D#���D������\���v�Ä������m^��`܉��r˟������܌H8� ����.�I�t��Tr"l�M���%%�lca�c�u̻2}a	���Jǎ�0�X�&�N��HJt��AU��|��@�/.�t�9�Y�!� �_�_mx0O:�j�T������33���6 �kYC�~i��T���{�@����]z 4˳r��fA4E*E¬����P�����I,ِP�Hِ����ϵ�|܂��a���D͖����͗φ�pT�	�!6m6��.S ;h�l�@(\����+�tE�i~='��e���~+܀�<i��3���M?+>��1/�� �4��?� 5��3i���J�^.�͖ydl������~��SokG�%���A�D�w�<$u�u�X3k��H�)�`Bh�v婩���Ⅺ�8a�K�_���`%$^65.,��`��]���-US����q�[YE��q�<��m߾���|_�O�+���/�*B}��X�;�~�A����U	��y�%/�T���Fo������`�ӎQ<��V8��f|GcaW���h>��J��X�
����>~	�,�NT���
x+�����B��(��<䦢������Т��#d��D¸D;��]���r\>��,���J�oˁ�O�S&��-���w P�mx���8�7��~�����W���c�흋����e� [B��ɗ��li���4��[����#&��0B1���kBS9��WE�)GJ�*
A��W��J�1�H&�O=X=�.����e��D�*�;XtN�W�3Y7Qz�P-�W^����̟�*�3�����x)�K�C�7��h�r�6Ȁ�lQ�j|n��V�{�R�߯y�x�2�m�JA&QM�Zs&�5��>6*�>P��:�uk�Ym1������ښ�-��Dh�����;�(%}�f��P.���+ ���_d2}�Ōև#�x��A�TY+���by�߄iz�����l7��*`3�����Q�C���^˘So�#�\��)/��'"��>�I��z�Q��<b`��&-Y(
��k��#���v~2�1��ctI��{�=���(y�3R�ʺ3\`�G*�< ��M���D��A#�Ee%ɤ[��/"'�������y0S�B�  �ג=@��:x��/�*��TGbq�����ЦP�70ni��,�z]���d@��-Ř���'�������m����y���ɺO��F��fGʵw���i��qX��/�@w`� x`�=���h!�&��KY��F��n��¤�M8\vv?]274"eg˼`�#��w/J#�K�����8����Z���ܨ�D28W�,X!�&��ӌ���|W����
o�@LR���]q�ᯙU�Ī��3�
7K��K�f�a�ɯVd����m����,���q�f�S�L�
w#XPd��*��A��n������'I���xч$~�u��h�ɺ�-X�u�l�EԜy� %\_v�oc0�:��{ӳh=��y4��DY���L"�$�*���R��r��[�}�F�߄�]ǫ��XnY͝��=8�9,#�C�N
r�6��j�ꄟ��eAQ��dd�%b חx��(���/-�%Mi�;�e��$:LWǜw�*��*���olXn-&e�`�MCL��ǚ~��-1�U
ct�p�b|!���H�yC�}d,�'M��<
C��sU��=
\�\$�����wGr��-;5\�����2i�<-)�If�B�oK��!�N�d�TTyh9�hn#�?�Ϝ3���,��S���L�u�m����6hj���τ�h�)��䛤�{>�'�y�x`�� ��ҕ�9����n� ���Ʋܬ,v��8I_m;_��.]��>�+xOb��ٞ�_J�� HӇ8cJ��Z�3����@'�)��~?cv%~ѐnz�����1q*�iE�p �.�4���|!$���"Y����9�Kv���Yq�k���� �]ȧ�8u�����S�*��T�$B�^'�P�ysE�+}��s����:ö
VY8Ro#���C��������&�_/�~@�\���EK59l<�����%[��8�� fv��Q�LWFZ�;�y��Eݚ�H{���J�ud�u�fS6�ui�+�0�}r 4���_V����S�)���Ve�ؕ�F�iN��܅f B[�}D�W�XgujU�=�LT���Wє��n{d���d����L$�����a�,G4y}[>�&�W���@އ�Úk�(�<N7�T��z��K�~gQ���b�N�Tp�0��C�g�${ܣ:% ̛�tcl�O`@1r9D_/T�=�ckia��1I]�l�@���:����^-�~{~�d�ARme���e�,�:����g��z!�
X�O��L�������6���:H��L�Q�l���D������
`�[
V3A�⪩�L]����ϫ�Tk�Q�ͨ���4;�j�>�	(ް4ׄpzSs0����.\�l�s��غ���`�Y����_�c�cr���K9�	c�n/P�}�5�?d������/��j�T��UKTJ�^�	����tm��ӄo�Ѐ3�}�||3��2��mfbN�~Y�7��h4'&o��X�7?��:�%�rr���خ���~�J�j@r�\�p��*�U���6Lc���e�g�Z���Nƅt� v��������T��l��gcL��!9R��v뇩u���(���D��M���ݿ8BE>�<{�#��G?�*��q��\ ��0	��]
n�$F���1rS$��h���'�c��J��s�9���7Ѫ:kI,Z=� �r�o,4�ZqUk�fZ�,��^j9uo	f�AQ��ь�'#�Z�]U���~���o�Px�Q3���:�!�O�9�?cO$B�Ꭲu��vؚ1}'w0�>��_�ˬ}�_�t	����Y�c��&�^|������j��Fu�C�[頉G���������&�0�K�9V���Gn_�V�[;/8��m�=��n���"��'��fE�*K���fOF�.��=ć���z�u�i��O9s����Փ�����I�^̽n�����,����OUѓ��/
u���0���{�,�=�l����tߥ�rt������t�Ց���*C�v���t�]�m��3�g�� ���x1L��
N!��O�r�
e�r�s�v:�̤�鏞Z.ˬTxaI��鑼R�(9ev�x(G��*���v� �ϒb�
�a��Y\�!���s�h;��^'IP.Ck��W���$��?Ōvu5)��\��U�n�g�fj����7N����3�J�+ǰ����p �|���y���@ŵ��R�v����&��. �q�B3���;L��@o-3�5m�#�z	vP���vXd�r���s��1$�k�m��A�	;�(1x��u�_����B��p�QH{(����rZm���������eO�ZߧOf�(엨�ƍ�?��O�B�D����ȵ�\�ɠ:$q��!�	��2R���R��|�� |n�;�û�D��{���Hzt�������6��<�� 1z(��}��r���ak�I"�%=�sp�jBg7�G3M��"wW_(��P�.�BH�V1�X\̱����F��ܡg��ç">��U�С!~oް�4%�����X�Pa6*�)tu5�-�y��ӑ�S�:O�w����sTh��-���Ti+1��oc�sR-��!�b��K��~s�����J���R���*���x�ɠj;�3i�,el���݀������:�i���_5�'��($�'a׶���#�ɧ[jl�Q����72bF����#|$���S�u�Q���d��	|h6����\{Q�O�JJ
v���U�����e�؞Ex���0��*7Z$��O��SxI -*��>��l?&�B�k!�y��j��9�!;��҄�� �d����DW�H͟}xs�]��L;]��L��#o
	�ά���K`򟚔�Z��G`�F� �ĻH:�J�x�
� K��|oq;�$��S� ��Ä&�6O�M��#�h�_�����0s\ �){5�$Jsǜ;lM�ޣi���y@M(/�Վh~���
l�	���StWZ̘�y���@�7\�����y1@M�n(dM�Dz#�v"w�H$]t1I��IR4�߭���[\��4�11^�y�Vh�:V��tI���mL5�0�y�� (+��ؿ��~�GCq�7���,�=�E�=^y�Uu����!K��[�RB^96,�w�NH�����$�b ��sc�W}�	]����/� ���i�g�ǓD�:�j�l����}�P��_��a�G�k�#���"��'�#J�\Ր8J��av͑L�A�O3���l�&�d����3�Kh�s�����Lu�L���� ��x��4�۔zV�D -3\mSC�����Alȱ���F�����k�<2:�W�w�`#@�rK� �9����'�+��>���iZ��~�5��ԧ�^rΆP��i"���4S��Β�� I����᭟�Ù��5�D��fY�hy��Ẃ�V`ח�����}L^@��H�⩍�j��FJ�z�S�jz2�EE����u�~�K�_m�մ2�i�%u��1���S��r����� W����S��o���6{F�/M59���hWY&���q�%h� �� ;<�_F-S#Ǘ&��͌�?p-`� �����(�Ux�ZD��B�8�G^�y�E�ĵs���#8�㹦�j���Ӷ��!���%C����p��m��D��Ig��QGF�*�x��S\����hDK�B��Ĭ-vů�uO=I�׌�Ŷ���H߿v�(0��I�C�)��axm�}d�>���:J_jh�[��� C}R�m��>�6���h�;�eC뻉OLO�WO{E_�K�fV��sd"j�W��C8(B����Š�/��?�<�D-���c9��fg�w,\;WL�.6�3�,g��E��F:p|"�4m��$-!^#���|�eP��߷;G�v.�/��\�!^������ v�Y���6'�J���a+���[�����h{xQ��{�f�&��tvMQ�Eivu=v��I�a�D��GB�����ߩ3�eZ`��8XY�m�+u��Z�=�Ǔu���۠�k!ŉED��0
x��w���Zs����G�ځ��*o�S�T�R,"TZ�n3uh@��(��%vOY��H�! �T��Q�-q�4��Y����OI�]�Ī	K���=���m��3�)tgFT �����H��/t��7�oc^�  �O�����_	>��rkz��R�i`w3��Gj��>����PU�:�q��\F-�T`���Nj�#�kJǙ��G�yk�r]��4�p�C=���ҼS��?mCU	�O��NΚ�wj"�#\�`�|u�D��/�<ɮ�R+����x(���+2������X�h� -F%���-��0*2��M��M�\
���Is��B�/�}.{EV7$�9�H��6e>h ��0�=׭_��}��v�W��;�?�#8;��w `��+]@�~W+����kh?t5S���b\���:�k���J��I�W�� �$}U���tIJ���� H�Aڟ���ŐPcu���B�_���Ԁ���9���� �~v:�5[��ẙ��o��1�,��F+�" �"�S�5��yݺ��P���<0�{�ȩ�x�|�ދ�b)"�C�;����U�f�Ni&N�ڂO8P��N'����~����e1�\n]E���- ��Ckn����� �?5� |2��DHa-.� �|���r��/0���������ZPG�p�l���h�`�r4%΍�ZYVB�'dy�|�����5F���?�"p%�} )z.Ur�"-F~ٗd�� �Y��V�*�L&��8�M��6���kzެ��k;l��J���_0�q�� �|gA��3>�9�u�4��@/W���;�3>�&�M�z j��`)93  ���A:��%�*�d~Mܒ�D� d�K1f�p�7���&�=b`���Ԡ#Ƀ�H���E{�!~�G�PLNi��f����ܨ`��lx��z�(�!Np�TRh�_�=vm�����S�0��hy%�EX���͔jʗJ�Ym�|�w,�s���`׵�R3(��� #5c7�e��d��v��h����RڿvrWV����/�<�o�֑�z��N9K�V����Ee�x�ܫ��ЫW�p���ָ�?}�͝h�9a�r�i�|&�@:*Py����=$����CmE�ܣO�!l�h�Z�t��G�.iD*{���S�(��/���b>żJ���B�`�����o�CS�h%1bحu����G-�j�<�/�[8	�iB��'s)���**�ĥ$G`�NA/�x]��.H��%�DzmO�"������Ӿ�$���G�6O���EL��o�\̖b������c��6{?���\zv:٣�9-%-l��Т��:'P3)
����w�<ޣ�.�w�c�Ѻڦ�����ED�����S�S��0ncL��zBC7/�e*{^��+	�ʑa�k$�E#::��E���{��	]�/�V��qvM�-q]����`���J�T���Ϻ�$��I���ѷ���8����Eʑ����"�)A�DT���d��"L��*�~>e���+:\=o�o>\sJ�P��-Wc���=�"�p���`G�L��|5-��*�틌�n*����$�d�D����M��W�����Ӣ�e���r'���c�����>x�����I ����.��G���&�4�,��1x�U�.w�J���W@2u�U+N��T�z ����[@�k^�1���� S�0��i*�'�B ��mK��b�Lq`�SN9�?�	;k)�ѻvRM�
�)an��&P�P�K�.��3+�R{��W�`���?L��Ç�#���s��3�
�V���_�-Qo�ޞ;�1�����tX�d5}L����p����6��h��]ϡw�-����a��[��Ҏ�A?�F�j^1v��%���$�?�/j!8��g���b�ʘ��/`Q^�B�)u|Lԋ�4)�����5��R!�߭d������0K4�K1�P�p����=�����/�0�(�O�u���XC����������,?g�mA<L��?���ܘ��o���9D��$�;�u�����L��X�B��2��%|�,�ja]1�(�Z����F��7[ߤhy^��V����\	���Mw �ޛ[7v�=���n�_y���Q��n�v������8uӬH�"��j���m�U��f]~GP��?���_������G�m�5��C�	�b�lS��D��}VM��2E��H�y�V�~�{1��A:N+���X�~���f��eӤyȷ�ڰ,(��bD�K�b~�Tp�*m��:���ɜ���
��\B�g#i}��6-q`Y��S�I�]�B���������u���:,f�o�au'�@�S �<�d`�j�l�!���|��N~����%�so«#��3���~�`�-��P�a�qO�&&���QC� �S�Ǩ<�#(���)�V��&!x�!���ގu��p�J�ɴ	C)���R� 깰������u7�KZ:��Ӳ�o��ȠB@_3$�����<y�E9�ITc�ː�)��O���0/|��i�e�7R3�W'f���ڲ/*Pn-�O�n9�
n�QS�"g��s����	b�]zt�-�ɻ�����ҭd��׈N��U�\ѻ�sk�1�id��"�)��CW�9UpC���Y�b[��
Ą��^�vh��d�����I����c9~��
����Td���a6�����
�����~�ἸBm?I�c��	�T(Ǒ�D�k|n��n�]F����Hp~�r��+�n�/�xWw�|������X���!m�\e�V,�<�2rS����I�q �0�uA�D�='Ղv�*8Ґ�'�q;jb*%�#0���9i�G#O��l�d�-1����t�5:($|h=QX$%��o��Ҵݓ�b�Lk$%F�E�z1�F��V�W�
���;�O���D�a0����<k�r"�A
����9��Q�VD�W��׫�����m^�������ƒ܉bܘ\~��pW�('�W��N�y2	��A�d?)��%�n�-p��=U1S�]�$u�אK \[��B��$ᄨU��3862Qc8~����Z6f)����䎪�&jJ�W �D��u��%/�Ł�pA%HUѴ��ܐ���d.���f�l�����x��15��_�V�>bE�����E�O|��b~E��!������vE-���v)��kP��<���A���6����Fz��3�H慠�ŻC�9�E>$5\{��dT��������,�nL����Ɂlp�>���)h�?�T��Ep�v���kN@a�q�zX,Mu-�|��@H�t����r��ng�l���Ӥ/�0`�R�s(��1���ח�&G�Y*�l!�Ď�Ty]ς���?0m����	�D������a�ڨ�A����Ǳ��	'立��"��_U�J��(}��2g� ��[�S=f�j���i�2"� �VO����e����=��Td_�e#�U�!m�4��<�_4��v% 3Yp���<��������to�v^�=\iBH��ٰ�����wKxJ����u�D�Q�Ȱ��g�|f���K�U�X�T��~�7���X��yW�:���LB�T����E�X*�Ϯ���sq��.hP��}p�F�Y������'����G)��R�x���?m�x{�g,�yC.TW���x�@�~�Z51���E�i;�C�<im���#b��{+�{����Q�l��~_8�`%�������)"5P/X|)��QI%]	y� ��?Z�MKy.;䒎�w��5�Ԫ�)�s��ݝ��S�����+�^��X>��QR{.���J�s�9�ʇ���@_,���}��X(48lO�T����%��u`G���6ɧ-B�����)�6]�(����x5�J��
$��t�X5��K���Kk�\4�w�|���ܡ�P�H}� B&V����2�ԇ�L+��6���{ }�ai��/-E(r��
Q��AϨ���}����_��T�/��M�U�N*�)^<�%�<q��qMy�����U��Q=�����ܔ���⥵����P(�I$n5e.I|7��oW�]�%>�>��L�{�cQ6����V3\	b`ٟ]I�ie,W���O6��B�X*LC�	V ����?�W[>!���=K��n�Q
#�[z	����Kk��N��b0����I6�����h�Jh������3��n�RlX<���hWKe��P�d��9
�5�ǉ��/����8jT��jM�2?J�&�������%�j�Q��n�i�`���8:�^;�<NV�޼�vd�yOy,n{��V�:�Dx��!� �(> �ӌ�w��l�F��P��c����vu�q�]ϑ�c�=�jޖ���k�3P�aR�	���'���<����s���������3V���	+Q�j��+�u.c�αF�a۪_! � sv�8���dA<_�ovB{�Bs6�o�������5�C��/*�#�����
�ʷ��
�����'�i8�%��O;G+<��n
<�ėj�m�=zҼ	s�A$Ԫ�(ww�F�;��D��x��&7d��z��W�ԎZ��6;����?~	8IcJ�vY�Y��+��̗p���]?�" �so�y�geI
�"zt��ԇ�^]����=�Ux��;�!�X<"(�(�ݼ�~j��WkL����S���K��R@�۶��(7�rI�}j/�$q����O�4pe�*�f#�@L����f>~t�\�
P�Lj�"c��C����Hh�V���nh�b��]�@��tm
T�d	U%ۋ�Rk����h�{�NUпͪVHGN"Yz;�}�tT�a������"�8l�W��ؖ�0zEҷy�p��̃���yY�(��5v�Y�E��q�0��F-�����>)q�߼po�g��	�.�aD;�4��_!uV�L_�ț��odb%�Ñ�~�_⣓���j�a.���Or"0�̈�b˕����. ��O(��[�O4G�Bb�o��u��G�X�8p�r�!��vŊ�u�_
�<�&����Z<G�+_v��9����H�C��ו\��NW� ���]2�H�<{���r�B�@�ʐ$,ֶxm��$>��Q��+�8͸�~S�h1������XOp�}s@���w{֖Un �����$w�����F?8&�#X����#�S�g�
��+S�Ќ�0������w��|��3V�o���jY��{�f�`�[����x�����2�N�~��7{�]HR!�d*���`��o#����h�@�V�4�.9����?#�̲MC�G���9W��(4*����,|u�tM�-4�_N7��)d�\Q��0ӻ�(���td���X7z	����V��!˩FPz���29.F�YwJI�<��n��ֹ{�Zd\B	���#�y��".)�?4�� ]E�pe9��]k-�c<<��	��Β��'����f_����6��,oh(�Ę멤�?���%:KU�]�]�A�a�=
��c׈4{��x���ꐤ��cJ��S�I����t#IBa��]�n�s?p����;�@L�,���ĩ���̖���5�S��L�dI�'��C���Ӟ�RH�S��r����b:�I�AL>I� ���l�h ݋��߯^���^��%"�<P%H��ʩ�͘����/�
��I�ݢ�*ŐoOǀ�v�s�~�]������yM��1	hZ����x}�j��
�-�s��X��^����5]�3�{������S�)B8��`9ƙ	1��\èڳ��,$����{������t�M3/��F��7��{h.̡�G�W C(pI����Ξ��dG ���Z� ˲�04��J�#q���J� O} (���:%D{?+��KE�&i:n��i��i"��B�������y͘�,Z������ET	�{�V���mM�	�����_fW��]s�6�5�w�q$1F:֎�Y�8�Z�5�U?��V0c̀�o�����[���VҾLBQ�j׶���Q����%�5b����|B$@ʣL���Ç�7:?��ß��I!�A<z�Qy�j-�"әpfr�}��N������tWq�o(�YV�J�$�v������yfN__�4�;�@�fb����p[��u�N��ԋ"J�g�vb�q-���tl�*�pnUO�y�pՑ�S��ҥ�X��z�m�^�%��A�-7�h++YG!� �!���\�vDh�]�	���BQ��T�{����0H�a"����Q��a�{�(�ܒ�z�z;�����vV�N�9�/'pad��X��_�c;!�K���GW��C�vNɁ�M<b��M�ia3 ��n��p�Ǔ�A�>������qI���b_:�B�&���X��W����;˰�cF�]��e���f��/U��6W&&����f���B�����
q��) �Z�!�i��p`�f�a��z"����&V����{�K��6�(��c�U�UT��)�!EY��G?=[���[ �ǖms���U������T��(ɼ0�T���:�3�-J��P{,�^g=_ߜ���i�f:�\E9��Xz�Ṙ�N*��l�h��Tqm�i��|!�>M���ylf��"�ql؈?�H���{�ozqNER5��>����`o��ɓ%{^�wWTz6�.��Q�d��t�h��M~D�)[��|k߽��m;���36�	���5i=��&i	�N/�W�8>�� ����yS4(��ב��HS�F�D����ȅ�@�W�+��<#Qb��ۥ��C�b䄀��p�N2R��4���d"�����V��e_�A�o�p�`��|�PךfJ�R6�����<��g��0կnx��d��|2���������*:B�Q�v%�R:/Պ�ؙb�5���ۖ�5EX>��A٥Y,K5;�JC�oA��@�^��Vv�j�k!TS��3���&m'\~�{������*��h�K��R6�v�P�y%���%i�%������u�+�E�4�x�M���xI��\I:��¬EHR�g3�Mu2�^b:�����߁��?\'N<�͑���U���n�tѱ�&	�CoX���@U&��B�N"��&�^�f�h75�LB��ylJ�޳٤��S� &�P��E��_ޠ j�/RIM��Cn.�������(|2��O[�l���Iڄ{�eb�FJu��}�wV��͖ujѕ�@f���ʎo*��9{^�͐qC@��lP
�Ù��n.��;��ș�2 �k?oX�N�{u������sYeD�?���`ҹ�{��Bf�#+ABR�^?�~(�RQ�8R'Յ���x�<��$h�^��������RN�0����#��� �U���4�2�'�������Y!��&8PEʄPt_e��K����o�]�I�;0ɗ��N�љaDn�B6��/��5Qs��\/D he$A[��IHС!��#��u�%�%&�^�	ƫ-K�a!�{�F����e�<uQ�G��7ӡ���N@���K���*�G��;�.Zo|��s,�|����j�)0��.�p��Zh�o�>x�8I�=� �0�1�;�� m1� ^���@y^ �qm�㥳�渤�a��2^ݧ��L\);"��>X%�m�j+�"#�u�8"o��>����rb���RT�cO�5k��	Vuv��	%x���	t��d�Σu3���6W��W\��.����<��Zb
w�x�Q~#�3B�q�n�:&���N�����de(���xP��,�y��K
�!��8�m,����m�(��J��9e�>��ё�����G�
�(�̕.�j�mC-����P"�3��'�1�B'=���ĸ�^�0��Yp��L'E�V����#���������[��̨�GPW��c9H�n���1�}#��ݓGu��X;�T��Q|�j���OSET��MU+ss4�� ��rx[�?�d��Z�,�Ő��٤`0��T.����b���;��e���>�{�fG�V@��M
&p�]%����:��Ŧ���-�� ���h��S�CJ�n3�!0P2xiY�Xb1z/����6�P[,T�L�%8nd��8a������>$1�;l�$I��DlE�So�=����j��&�?]��s
�u�2��m�ur��cTy�!��&�/���������$u������"~ɦ�H����&Y�K���S�䇜r_����Rrf65��-?����=��q�֠E�dc�T8���Dcu,M�	�n�T�5R#$a �����Np���-5
�\�Te�#�Tpv���Y'���W���Ne'�/0LUe��#�D���K��n���ݵ�XS��Z	�j��%H��N�����Đ�2��Yˆ_>�e�D�d�&FF^9��%�Yl� �t�l>1�>k�h��ʃ^���9��	M ɼ�Q?��y�/u�n^���G�B.���?t,��͓:Lx`k��L��ܹW�ͅ����J����s��:.hmAۘG}XF~�[�l�$I ��l*�'�r
BJϽy�:?�_zzS}�~�YIQ��{����t��Z�y:.
�8rA�k��(5n>B�)�G}8	�_�H�S2ّ
<iƜj���F��h��&MaO�:O�Z_^?�����-�8�z�J�=҃~ڈ�,#�b�����Y)�j �[�44M�R�t�Qv�5��eC�� 3#���Yhee0��=�_. ��7&�FZ��l�@������Ü��)�l���,I5�r���`����@)���t_k�x\���}N��}o�X����e�4��(�����`�1�t�*�ɁEX���vo����J��T�?�]� ��*/1�q��h7+0D��Ip�%�ɳY"!r�	��1���\�D0�rY���qX��%w䓄ƮPi�����N�� Z߰P�<3�yO��1��i���Ax�l]��<Z��W���2@�CY�c%�T�ө��C�>���%�`�cb�v:�����*ݤ���v�ԉ�8Ѐ�N��N��@G�~����,�ME�]U��_{fPr"x�(L�n�7���,i���n��K9@�"�T���wLh�@3��\�hx	��yq�1C�=DjBi2�On��w$��u��#;�P9�o�ypA��7�E���E�h�wX@Pp���*�559D�xQ39�VX�����p+�K
z��%�sc�ƕj\���)bB�� � T������yk8�o�'P��p<>��u�V�E�{
A2�N���r�
)\��Z�@�S-���Ih���oI��i涶L,�V�h`�jŴ���w2]@�NJT�$�;��p1 �[a/������̡_!�򽌫�@�4.B#� �,��EwbӤ�*D�L�����Ӝ����v�t����_��#\!�OwN��̗D5dj��1J������)r#(�2�Յ��]A����������U�W���">w������>�l&���q~�"�4�X�\Lv=H�ǐ�Z�i�K��F�o^rN��*Ѿ\�Hc\oaX�Kg��.���͵�t����0���&i��������3��ֹ�e���U�!X�]D�P`t~sN�3���f��b��:Qy���ק�x|��U�ѓ���i��N�"���ܑ�Y%�'q"$]#4fn��,����7����;
��|�]�'��E�Y�~��O�K}�/!�FXL�dE�x����}��������}C��1��=��\�T̀8嵝���   4Õ򏶳�g�e���."����w���h �����4�jguu:�h���I,�Yn��K���R�/?��&������3��1�MQ�٢�o�+1`��|ޏ��b��|F�BRD�sbP8�7B.��Fw���������U"d��Y��k���V������L��f�����$أ`�s�w`6�f:�&�4���>����ԔẎ0�Ѓ�$MA�f��T�!u'�r�"�����X{����-��	��G鬅��|�$r�)��n�1�G���P��;��E̬����/�l1(s�?�:/]������,k�)�qq�~� rdM�˲�f�,>D,�kP%o����^��d��\���B"�]����u����S�/�"�j��Ŕ��x��/���u�q��pK���U
���&?&��x%�h^Rf�:!�2L����s�h��_%��7+��`wVҤ'�0g?I
,Ww��B�ºt��K�_I%s���_4��c{t�@OlZ�G1љ�>�,w����G]嵼���ٜ=�ShU��N#�dš𩘠�Ŝ���a�Yd�-6]
�ef6�t���(����_�)�ɍ0\ن^�o���j�ds��a%KOb�e��_J;�萶����/2W�����Aێ�ie%C���:;��I���Ǧ��oA\3lc�POu>HGųy����Z�� ['%����*���<o�^�Ɏh���;�J�j(��Lʪ��ɓ��A$��ur��i5������bhw/�%/�e'D)�O�kP~��.hK�,	�s�ɲͧ8�:�T-�M�b��O�
�%ה�y�d�~י����,/�g?�{��B0��\H�	%�Ue��
�ZY�^��	Ub!Y�nV~���~+��:�/4�w�ݰ��k��E�Q#����mhf�d�ݻ!Y�>4��o��h�/o��l� � �.556(�s��fH�. �h�/}�K�7�;���??�jn�Wϋh����UЏ�~(�W;�M�y�|Ylٴ�}Q���A�6����wg2����9�j��l����fr�G������3��h0w4�ꐊt�5�8X�?�aGc�j���ddk�:�o&^� ှn�zG�������Z@Y�=3w������t&Iws<
���X��M�0��5�� ������'�a��{�vq����J���an������u�5Ȗ q>S$�G�aR��dS=��n����2<�t� ����`�W5����g*�$�%OGJt�c��B�t0������k��WN�]���5 ߿hw䄼V�15��$���n-DϮ�E	��Gᲀ�R��_I�%�4!Чkc9�H"__����B����-e�������g�I��t������Z�\�-�8gce��B��&*��j���
l]�������~�����_����H�%����p�ؑ`5����p��W�Ќ��=[�H��T:ˊ�.#�o�K�*�W�R�%^����s��V
-p��p����]k���=�y�0�V�T#.�|��-���V��e`#��ͩd/���^�;�n	��]�v�:��ˁ�G�½(�Ft���*1��L݂����3�MR�oQ݇�qs@�Ͱ�g�>��?,V~�2 K
��P��`�ߚgl���*�>/D�e�wB1? t�<^b������4�{\��<��2�(�}TtH��n��̭ �2~�����q=~)8 Ń<�Q�.��f`��!�T?���E@�VJe��x��S�ؤ�>���"wQ����wT����(��3"�:N�r�Nq�^������6��Y��@�3�T�|/��Gtsrz�"ႻS�5�@�x�����|T����%�x4ḙ�����fa�7 �;����ً�Q��Ϯ� �d�sjRv�WT5f���H���u��#����8�֝���2X�ٟ&�����g��`�P��-h��F7�@��k9 WLx�aߟ�ۢ�?/-0A���H*���|]SBS�:f�]��o��L0kp�N��8�S������uY��h,�,а�8�´�o���ŷ�@���Ǩ���jCT��b�+�E��w���T{ٸ��ˡ�5�m�n�����\�A�ǴuM�w�}yq_�W�
��t},�&��)wۂ�1����w�����Y�w�����;ү6z���i� mD���l����D[vy�g�ۤe�>y�/�5K��E҉�B#Bck`��ު�0�D��bN���eT�e)������7�|A�|�5�ٻ
*�jI���B'��bܧ��+��zȄ�n���� fX(\�����������Eߵ��:��hX��Ou�s���V2gɊIZ�q��U���-1̶2�9���~�r�)Ѩ�&���I,�e���ZV2V�ˠP�ϖ[8\59z،��,�א��	�&Bk� ��&>��.M��J�B	@2��Bw5�JR	����We.���,����d����!V���u��Q��y��-}����ڡ?��c� �{n����#�S�lw�vn�B%�Z���^�o4)y��)����r!�g�����5C>ȑ�O4���.��vp�=o'��ׅ��3�<�aE�����*cZ��9���L�� �A�}L���X�w��3��M�g��M�ѹ�@m|C1t�� Aه&X�aC	���1Rɜ"�	A}�eဠ�P�T�y���1��7�.F�i]�]�Y��;��-a��9W60_x��2�"y���8���^}�y5��]��~�!,�vi$�;�p�#�b��uS,��8i�m��in�):&k?X0�ۃ))���L���CFW�b�\
=T����m�8:h�o@H�D�U�����[�hYu�ֹq��0+�]�1a�:��98�A�����(e#�����u�0��1�3j�,)Oj�^Y�|M_��bZ�/�d��,���Wo�������e��Bb�.@���"?���;A>rkX�4����!�ޘ���j��Z�Z䰰.�otX�`Xd��¶�Y���ANV���kΝ���.ސ�n�z�"@�4Q;c�z��-*�^��OH&vr�%u!��{�!�|�[���2%,u<��:C��g����0�0�8;�tG�\@�0���\������Pd�Y^֧N��EE�F!k�\�GR�}�?������Cy��L,�,}�N|�8來'z�Ȉ��.eڗ�t�.�H��6���������j�w[�s������/���Z{��#��W0J�s���2�.�_m8Ir�7灴�rp���Lzwj�-V��<e�:�v���!�E�,X�W�s ��n>  �]i�*I���v� `^(�M�8���Gf,�X!��/i��p���֍i鳤]Vb��A�x8�7|~������W4�$���F(ymk�����B?�(�j�X��V��R�?��ӳ�?5ԂT��l"����ed�bz���!�kh�kP��$=�*df!5,�=�^P�
���uM\5=�u�����<K�4Љ�����h��E�P)�n#�w�9��b�ЯgZ>�)�<�x	�;�k	����y����\���Ձ���Fk��M���ǵ����q� ��U��wNR���z��;~^L��7�\�SZ�K�ڒ0P� &�CO��oy��TzƉ����c���4q4Ǌ��1S��b��x�X=X�� ��y�A��,�X S ΓR�7!��� ��<�R���m [5i��K�����*�rBy�k`ǲ�B�:�`b��`�D�۵>|�'��4�Ȼ,�\���ߗ=�YL������t��	qM�F�F�"�,��awp�@bp?�y�9q�qJ�(�f�Q�Ǒ�N�Rs郺�s�<��������V���w1N�r�)���n��֐����U��2��ձ�ݐLb/�Fګ�fDr'��ƾ%�""F3�X8Ǥ��M	�?�8��Yܵ���d��G�\rR�dlf��P$��0g��tPs�	�^���;���H����/����6�;RO�/)+t���ً���5�EĚ�����%~�M�yG<Zm�	~�e� ~�~K٦{7�v�d"��R�c�"�7'd�O�S���*�`�3��1���:�$
ghɪ84B{3JO"G�x��/sc�>ݐ��3�HD��=p���:YR������O���W�0�|�y}s�x���&)"3�â�,nH>`7�!6���3X��[_�R�����聿lc��j'h@z����;�UG��r^�S�(��5$�x���	��xCL��3\�����^P��p���E�T��0�_|��о(C��.M�i*r,���>N"+~��^.��S,�ocC��ǫ@1��W�2���Me�9<�8y�6=��G,}G�d �3�+i�.��AC敏�҈s�P��"�I&C$_�b3���:=�9b��kߟ��m-�Yԫ�d`�BM�0��܃�����B�=1���"�te�S�X7:U7�M⾺o�x�W5K+K�:��{u������� {�~֖�r[��hn����(-O���ʛ�ͮCB$C��y���F��%�+�u�K����ݢ�R�j���wQ*��G�nى�u�vF�����zDR��c;�8� F�7��;>�:�F[��Y�-e����,(g��VRڇ%�΢��7���{Z�\�<��?���+LE��H�4�5ޙ��<��]��M�7��8���f�����^�3*��j�������o�O2�>���biF�K�?N��r�ԠX��J���AN��O��SԖ��;�k�V�J���0P���o��_���ۗsb��f9dG$D��X�dQ���j8B��]�i��ޝ(�g��ʠj;���R4G���z��q/�;$C�w�-!��gr�'���}�#\�aݎ�nL�9�q���'{AZ�Ti���]�7�5��VL�>�����7��y2�������[z%�/��J�:02�~�t����Pv�9�T-�X�H� :-x�������c�dK�*�Qe.����O'��d��%9) Z��AK��P�h�-�V��1����w�g�!�%̀�P
��!kV���ŊjX����
�����Oqs�d���9Z���TA٦��Y�|
�Q��.��K����sl�Ds��h�ul�i@M�s^j���ȶB�r����nCcl�B�l�Fe!�'���:��oL�/��`����)�����L���D��RwT��/�J��֏�UI�父:3�#J�m���}=Q��G����ln�]�<�1�F�����ͅ��hW�4��~���v�.?谲g`��+�w������Ӵ��~�9��x��$��)]j��B�;ow�[ߜI�|^��/&�b=�y��>݌	����O���\C��/�'��1)\�`�r%>�4c�=�$!�}�3�H���	�Z �������S4��1�۷n ���&pV�I�����AŚ�\��0uD��R���~���ٿ ��!�!��|�ZyBwV0f�r��D�����e9b��͝ģlw�=�"��(��k��o3���:���,c��i�,��R@������*�A�+j-j`�F4���T�"�P����z�@�	�V޲��6�Koy���e�V��-�GX�m_�msBR!z��\u�~�t# ��T���7w����Z��h���Xs!�^�e�?��-ۻ���Άj�.�șJ��s��m�h��!$0�W�FOx�A\�<�,$��5�G�ݰ��e���)+�\�&�0bniF�:�WÃ���X��r}��
NV�	rİ���N��&����ݮ�<�N��^��_��Y��g$)%��(!�hR���d:��GŴ�9���WM,T����K�5�>VЩ��R>[Ģ���U�����CL�ǹ�A�|��AY-�maf�l[uj87���H���'�#I���/¦�3�1�T�:K	��B��PAʲѡh_��p����_�{.@�A�����<��Ϋ�>��dj0�r�΀>��0K))=_����ȵ��`��M	���]�1�3�F��y+�ar����x$�*p�E��)�[����f�+�*@�}ן9���|����yE�ysX�9������)ne�Q�HxpjWP7�T��-R�aW-�M�i"�^w�8�dn�l�im�)���C�0Q5����r��T��WC����P���)�މ��#��m\��B�{���s����i���A��*�����1`[��D�e���WY����H�Rei�aJ����|���'@�c@L#��	�+^�l_1k��;	�$�V ��f���� �Igyn�>��� ��9�f�E��4�����pd��U��(��������a���{�i�W�o,P�����K7�-B!��f��'�. 9+����=�'�a�\g>O��Z�����>^b����1Zܢ:7f$�xٍS�m�
�ppϟ�;"����� z�>������M�f��IC���'p�ld�����>���_�X�=�����I���f	��0���Q��v����?7�2���q+�4�;Cc��H
�)�k6WaC&��'�٠.ԺlŮR&�E��u�=��1��2W-0����k��8��\�:a;V~��DG-��u�#R?"b���~p?f!�S�L�*\2ӵ�����n~d<��P�vˡ�?��Jz�Dc��a%�v&��[�ڀ4ժ�.p��'�{V�*f�Y�^�]��3x�5
F�F�tc����P7� �Rĕ�
����|��c�ޗ_95z�ɯ��q��B	q�9���u?�j^m[�����k&0���iE�J=9!WD�dmV��c�c����|��/���v�ߥ���T���8�lo�BK�v���p�:z��b`�/_A�\{ɽ��X��R0��^���٭.�LPo�5�F ��Sa[GX.t��;EV���Z���7N�찰	.����I�^��7����M����Tݺ���&9?��CK�֧���&(�Sl��6���H6�Y&b�sA�,Jg��y۪���(�GP���uO�|V�k�Q�a@=���� �(�܉�:��\g2��]_ʙ�fC仱��W��x:�F���� �j�b���@9롭��n[�1���
�l^<���5�D� �S�Mxc}����1I>r�9E�0�d${z��?�HU��mUp�8��<��A�|Њ�̔�Nq~H��mC�Q�5��be'�d7TDe�}��MI���2d��O�V�ˍ]}���~��r�El1k'��@=��W_���J
��;[6��9,�??�W�N�����A3�x4����"SĽ@1}*ۉ�㋳�&��Z�0�J杵SP�Z�oS�"���o<xc�ؗ����@4�~�}=�q�Z�7���B�f�ަ$��n�(���4D��D�`�rt�<i�ǱᗷYˈ���8k��yX������#p�b������T�lܷ/�╱��>�^đk@7��K�������N��[�\Pp��汿�$��v���q�a׬������"�DbpI{�V�����,5�:�iM�^�$W�+%��B�Q�6S�����W9���ɜ�O+�J"4�?���Ǉ�hR�1�z��@��L�L�=O���m��(~?�F{�O�٘�#��+��J��Z��e������c�e�Q��^�r���al*wd]<���a�ͭro4�����|ʟPB5�������\��%���Գ�O���ܒ5ߌ�K>f����_�L���_�� ���壭�4��Ύ�Z��K�:���"Ӕ}FM��������)v�N�Yˋ��ۘ��w2�	�Bc'm�Ȧ��D
꿬��}��7�[����S��!�V�U��N~I&Q�YWW+A?����"�}����<c�]?c����/�-�'�X�D�Μ�+a�;��X�R\��h�o��ְ��{���Z��H?���/��Ҿ�rc�o2S(^Ν��5�C�?3FU�5�g��~7ӕjyW ��:�j�j+��Md� - �mr����w5Em�U��2`�4�gQ�df"}�Uw�aW�Eí�%�σ����
UOj�!��Y������7i����Un���0Û�W���2�������.�)os����ѹ`���g�m?
<Kr� ��Q��Pq"�R�e�	4>��=�u��Oa�Bv���A�F�ab�d����K�)�q��t�"���3,���\�xI��a����2NI�v�p�~��6���3���.�a�}��fK�MՏ�n�yѦ �n%����L�<2��ڦ���w���tP��ͨ��*��E�ٹ�S`M�P�^&���B����[?5F�^p���L�)�̌7ԟ�K,����;k>P?����ϓ3�U�`1V�?�yA��bߖ�o�-���.�Qs�SG�;��8g�l�h��w�rd�M�
�oLC�	n*�"�!{a��,$�ȟ���%�T�4�N�S�q8��W캬��I�5�B�#�z@W<���&��!II��틅�˜��v���!�	�;��&�w�Y���i	K%���28�� ���?�O�
�U:�+tq�}!pl:B1Vҡ��ۇ�k~v��)?��3�I����7�Q�<,h_�XJ֞˓����#��� ��\M�j������\?��-z�-n�ι����2��/w��EVK4Z�V	Wҁ�tBi��^W�����K��DJ �����Ϭ�7���=y�tV���;&m�y�H��G$X!jR��NMjD�׋��c��6O���'���nj�7���|��f�j�2h���&qҐ�)����2{rV%�=C	)|�M�l
Q��7�a�@t'��{{|Tb��*b�e9@��I�&έ�`M��Q�qJo��Z�q��]��x~�0���Ͱ>�ջ:�p7�>�/�d��C��\p�������f���:��~^��s��j��R�?��X�h�xl�!��ۭ6����y�e9�-K�b���=�b�k^�[�V�|0�7���B�C���!X���
��,�
�sΜ0��r����G�914;�t�k�� 
o��\&/�i�B�U�m�,���8��] I�)jQ+���L[$���'O/��z�#�&pq�<{د�A�"91�Fˑ�|��L�v�}��f���W\��mv��h�Jz�ɱ0=%D��Ԙ>���E���O�Q�e{v�*_`��ׅ��-��=R��u��͞����ޏ{X����>̦`'9���$�����9>X�`;��z�y���\�g��� Zd�bW�L���M�^[�*M�l��"7l@J/cp/ɣ��T	; =�)f�dHx�"��¢�P՘���,hci��ҎLv.m_��poXH��*��zg8u���m��-mas��l��϶�x<���8������ָj�����,+j�z�k�+���ةn-��
����(aL�W���L(@[3��9�����:�m����ne�N�k���\V�Un�u٘P�J׋2��"��YrB�Y����S1�B�ʻ�����J寺r���Z<����w� %Y$+|�K1&t���	�;�y�HG��]���K� �ځ��)�i�Ac%�?� ���f ���W�u�k%�9q ���\!]$���X���+V��1�.����������O�H�z�̇bG�S�QBim�E~�&�}?��q��Xf|t�F�����%�N$�b,�߈�����HK�U$����򋄊�Oq�q�.O�,Ѕ�_����]q�*�����d9�h~�'��e+Ǥ����/@�e�.�+ �!�k<-����5�p	��H����c���l����L��wœC����b�k~D�
9��{���5���k�=��D^����u"9�/��%N��n��lQK���"v��C��[�GT)�|C��c�A5�
�0Ǖ
��	���M"�kn��e.��if/!�ş�:F۪�L�vu��*R��4h>�rb�c1͖�tǳ��ޮ
��!~K!2�k�,�V��R�Bҷ�9(ܸެ"+^�ρ�Te��,��Qf��k1TK���B�J�Og������6�1�eq� b=m�'��|��� �c��B"�NO���D�khY�ݹ�ڙK�#�j���3�e�G=Y��sJ�.��i���A��jN%�ã�)�y��&S�6C��A�N9yd�~7�DPôD�c���8I�!�]ز7��sN~"H��u�t�چ�Y���}E�u�Լ"��,�h;pO�����د��A�!3��z����\R� �p�#�A�*����&��r���"=�'֍4z*
���H��ag��MB���6,�uL�Eay����5p�0	8��S�k�O�P�2s��4��y�&�qq����=Pc@�mCv^D��0��C�j��!U3�gm�86�\�e��\cq��l�Hԙ
�^��&˵�)��l���^�'x�԰iT4�����ûl���_�V"Q*����@�f���8;�����@"�u�sE���S�W�ˌ�!��;R���2}Iy�>O����J���}�N�:ݨ��~�mW���p��qt0O(��i��op`uV�Q��H)�3�݉%�Hz��+*�>�G��ؐlc��x�ӱM�4�N�
���Iv��E
��|���2�B��!�0��r��@���/�W��U�����f��-�z�_��1V�cIz�;D����1k��Y-tt��K�T]�⪂�D�^}Z��Ց_۾�W��S�7�Fa�|7��(�m��?c;�8��[����F}�+I\2�|G�`D�t_��*�0�$���Po4���/Y��IB���7UnX��9{��gH?mA�A
	��	��0�9�����0�������`���������4����Ki{5�,��X�;\{������������ p�A���Lp��E��|K�39!�����L�����d<���)~A��d�+�Wֆ���T���6����_Nː�dJ=��/����� ��nGg���92�L���Ȫ�$qm�Vh O�}�&��;h��k:�5�C�ێ�J$��:�. �+օ��1����g1q�Q��C�c��{�@�a����}����*-i ��v���݆� +-!�7�wܺ����� M�Y'�LZm�0h���<��Zʛ5�s��"٘	��M^8R�<�& ��NT8�H�ou�j����͛s����]�*��|LI�^��V��0cs.F�a��BϢ�[���2�z����[����T�)s>f���[����0����8�I"���x�����r��$�.����v�#hL���7rli�ڪM�����G*8�$�mW6�\b���2�Y�b��6�K<���G
j�v8��ٓC��@R� >,��Y�WtI�xّ�B���k���p��P`O�(<�	�*�!U�Jl�ńR�+a���p�I+ ���Oͅ�!sZ����:x�p6�^�����-P�H�,��m(?�m-na`�"���d:2�Træ���#�،{��$J�!X�~l���kv˘�l��'��]ɝ�L1V	����
Q���aI�C��͙45�������W7"��xn?y��r��0�1v�Ph1��U�L:�b���҂ ���פ<�!�)�o~a�=�`����M�I9m��b�l����.����,Z��aQH��j={�y����2�c�q铄�� �`��������iY*�����w2��  ���2U0��}4z�[-�p-xl���9�b��t�<�*q��,ܔC�FaΖ�m t;���>ېP��8{K�Q�o���#�|x(N�c$�91G�#����zl��D|b�w�tN���)d�*�[�t�ߏ�|OF��qױ!p�`�g��)�m�W�����`��3U�Yh8��s��C��f&F��64~UhE�{'�_ݮ��k��W`�/!1�"�ݲ�L�!;�hlg}��LO�F����'v˻Ԅ�c?�0��a'~��ƍ7�(M�l/:N�y�O�_fHy�H�t��,�c]�/?�:�-rv�4$]� L$]�艶����:cv�#��䞋Re�������T�Sp����7�s��/D�h��V��U�9��"Xl������tx;k��n ����Cj��9�-僋�	��c�2�`�1D��O!eF`1����2յ\}'ekv�Ⱦ!�]�C;�(̋�?�?9eI9��+H��`x��D2�A��6S�aL��C�Uo
s��'�4XcI��c Y��'�bD�G9gEk�_Fm2�q�.�h
o�\��,b��� ιi�y� ��M��{_����lEq�2���G<$�#,��J�69S�<�}fw��T��eG����~�ZG��0&�B���b{�C�Y���b�ிM`�_r��Ld�0g��$��gZ�m�3BX�A��D��Ǝ"�d	��3:���0Hu��Q>ci�@�Qs��'Q.���-ޙ����k�Jv�{ǰV�����s(#�d+�^�pa-�@3|�w(v���=��#?e݂�1S^�}:��4�r%�'�����o���띮���/7[��Z�	�zg�s��%7��!� ���E��Xy��&#�G�{��`��s�\$Ш�=���{il�ti�������_��=��;l��8�jZoϱ㚛%��Z�tnm��Ɋ�h�;e ͙�I��qs�R��׾a�G*�Sƙ����,�U��,}�;�~M��z���U��g^!P雺uk�s!��'���ꇓY�z7���a:��#rjKN�<�9T�+�vc�t��-�����_~g[������J�=[~�2V��d���6����!�]f�]��;��īUe��eQU�l��� 7���W��$�y�\	�F����Cu������DKʎ砃��u)|�j�Ru��G��_�$�3��<���8f�W���������e:� $�w9.ߔ��zm\bV&�A���ޒ���v���i^����h��j{�O�(k���;e@jIUYL^!C��ڼ�ϵ����6�a�#bQ>�/�E��4je���}�㮙W�I�-��i�&՝���㶖��=�\���)�.<��Yg�u�Z�2���$����!mN9�P^~D#A�UU�%SD�ٲyc�0� �d���v
1E@�:�(��H���7��ĴO,�ν�3ck&����/���\V(�G(�L�# �3����v���L6-�0��"�!�
,���Z���MU""����.3su�i�4S5s��(CK���tY�aE%�VM����(B\!�R��E��;��َ�YRu�����
���!�`�I f��^��,�y%����'Án����Z�s&�D�v��5-�T��$��@2h���z�/ߩ��{���D��.;�ă�D�i�k��?,cT��jFc�<MS�46�O'�O$��S�5i�d�0�����{G����2==q�_�JI%Z�&�G�-�^V���lHp��\7�8!��s2�P�B�Ǐ�n&���n�6Um_ĉ @�����*���siP��Z�Y�E��`+>ÿ����=>"�
8���R�g�/I>��1`��O����}k��'pn�HK�Mx�BP�
��x���FW�V�������>dFFz��j' !�R��B�Y��KC�qm�sa+}�;P��~�_{c(��4O��.m8JbHO"�T*�ӠpV��erq
Љ��}>{pGG�(b ^�o{�Ѱk����Z�g��ȣm6yf���*%������c�s ��D�"<R-��,˅Y�vs7�D/ʌ;���T�7�5[N�(�!��6�;}��H&ZW`�?��cD�dt&���3ޜ��^6�^R��W�%�*�*\	���$a����y�)�%� }'��	�nx#�zs�G�_��O���ɧ��@�#c=VW�/�"ʱ�ow�g��k��!��^H�|ǔ7�8t��8�����K�Q>��<�u�"��*[�K�p�ҍ���f>�`H�x��"�~���¨G��K2yӺ����zt�v���C+S-U�92�Ƨ�/1E�$�D��{���s�v�Uq�O��R/�R�8M�㬵d7-"��B���W�h��"�8H3��q���o]���"��"��L6�`�3{Q}��Y��ՎsL$�P���T1�jcS�E���Z+�Y$ŧ��T(2��&��C,\���\}��Pa)��Hfm��?��9K+�.="ŭ�l!Z-��G���hR�]���$SATCD/T���6"�0!�sƟ](�h�j;��'6\�2@.=!fkNX -qkW.��o����M���	m�2g�Cy��
A66�A��n�g{��d��*�)u*T �*���}Ț����?k.�b�7�n�����H^VUe���,5-�$Bf������#����{}z����^� ㏉Eq�����.�I����^7/G3��-x^1?8�1�F���|=�_�r<S��q�P� ��DV	���m[�j��
5���>]��R��ɦ��O�E���L`��J��f�ڰ�����!'�#�Xx]��D׿���ԡj��p�$]�
�!,��w��'�6nT�8쪌�ؒ����c��9�w���fx�k���p�VӪ�9�%R��z�?Ѭ��BE��ƿ�����6�a��ʃ�ҫZBo�;��)h�����ծ~L���D��|���ߪ�_���T,�k�/�t
3r����^����Gj�'�ӳ�{�*8��zO�b�Q�eb+���Yu,&-�8�-�"T�{s�u�ڏ酹
�����h��|����4ǰ�ƃ91��6[}5Ȋ�.5+~8�ԍH�Yt�I��o��+B�S�(���ӳ��j�f�K��������R*o4,g�>�Q��0zWi^[fP��T>T#M�@_�f���y�ʣ28L�r\�/.�袽�e�;�����Hv5٥r�冗��1��G�Q������LGW݄��n]v�|U-0^t_���3
�M����2Z��1��踪x�8��UK)�D��6��� �:��#��v�FŉҖ����d��|�?ɠ'�5����0T�!)x$g$;Q�m���ym����y�;ufx9lǢz��j�3��rK�lrC`![��ъIIS�������_��y7E6���*i�>d�Tܜ�҂�!����R�ߧ�v���Z�W���j��� ������1YrG<��gyr]N�����2՞#�9���'�	�S�e�Q�	)�U2.��V�q�S0��t���T���V�]�/U�v�� �[�����2~˾�ZB)*�.�l=��{ӡ��r�e�<3�0�J�������(���jCm���$����$���JM����X�݊�EHU������o��^@��n�hq19����n츠�M�?\t�k����+xe�\[��M�1D2�LP�� x�V�A�|�����P�u�� I�-n4Z��#�	���[�QG�3q&^tR��Š�o*�H;T�;z���JA�d�_�k1$�PR<g�c��1U�3�Qq�2V�����ai����li����V'���q�]��BHZ�V�N�oixT'?�M�6�����t�=�;�Z���70
��������d8���Xu�?�n5-��+*�9qُ��Q
h6KOn(s{k�X{�����MD
��I,�b:&G��m�����F�&���YDb�P/"$Ecԣr������gڿ~�,�����
2��^���>�Fd7r���̈���sέ�Y;���o͐;!�����`�d�ǬƝ$:�Co��C�!94��s���=��K�j`��l=�Ut���>������2d��.p�W
9�(h�e]GM_��<Thj�u���ϨN�\H����� ?�d:��ٽ�9'���fn�'6�i��FId�146�+vf�9���I%�ۡ.�/�)���&��9Q\�g��B����T7f���a��[�/3�^�K�� ֊�5���N{�9���8]*1�@�D����-'���9yp�_#�f�0�A�gö[�DK����+���	���.�s'C�[{P�`.�WT����u	�|������0�.O�C.N�"pC���CoxB5K�TH�w;H��D�n����K�U����Gϓ���?�2 ����	H˰m����V�����Q��S$/�\p��c̶E�t�>6��|،Y�P���AZ��ho�9�l�/�?���ۺ���ZY؁��M��y|���<�u���a�'��x۪��U&���ky�}a�o�c|	$����PZTd�^Ѭ��c)1��%F�������:��⬙_����'��;m^9�.f�$�L7R������S9K�tͺ�	�b��5t	��pZ�a�)��>���!�/��ٓ�hcNw�5T�L�>ڴM!҉+�-	���na*���/�;L`O�5�������x���c��/�[�:��s�^)��[��?�k�p�b��������8Y�MJ��d߿��=���;�Ұ�j���oHXB�^�0E��6
�ݰ��30�8��W�Ld��D�� 87����1z�EY'v�3F��f(|ߠ�M:��׹�xɅ�i4*�Uvv%f���e�{�K���*���Ɇ�i{ɛF�D/mNZ�yM#�C�&�Yˣ��%�C�8|��HN�1>��\�j�2H;����܋�n�	n�b���
������Wƨ��/�����5H�9~�|q���Bv��z �)��1\�(�)�.h�gҌ'=���Kr�g��u�#*\nU^��)��u,`���Dg�K����\�ǻ:���l:LҮ�ׄp���p����РP0�3ڟ����X���h��Y���%�^5�ő��g5lF���Y���!�(7;�z{c�A(z�y(������S0=[!0?�,����W�8t�;4�H�&��E�2�P�5��n0�v�ۛ6ha�l��8z��c���e�(����S۳`}Tk�a��'�E���.�W�8$�4����=<нtٹ�~f�ɫԈ�vE�c�	*Og?��1�J����u�MB��G�.�7�9ǳ��<������j�8�ؼ�~f����.����
�ݺ�%��ψK��p�	��ƒ�	�}O P���z��&M�"��x<��3#���T;��D��znMm��a�Ї�h���׃坘A����m˥��SM�P��LB��cľ��젼f�Y��Ə��ik=���O��#�8�0����Sa���D'�|}�7)�s��Ð!"���h���P7�	-#��`йL���oG/���4[���cp�j�+�9W.����d�\QJ�g�.j}ޤi]w�Y�/�RB�b4ƑT���%����;�Q����i���w&�-��\��� ��(rlK������L�E���l"�3e���_���
��C������&[�VX2�:m��랄!�R���cAG�+�E֕zC0=jsf5.���h���|J��:w�Q�<�Ns���S�Q��:��:wm�nN^��7Y�ыʌS�_����y��z�AS�Oc�[������+2��a�쩐��UE�&�=�߱oA9XiY��h�$䘹�]P9�,/����6^�X/v�{C��\?���p×�խ,�4w�F����fo����G��=���JG������k��-� '��1��O�����7k6��\M@�Ь�� m�p�gg�:9ּ�@�h��5 O�-eD�W0���a��]R&�є�1��kءM�ҭ�hc�V+B���_D�4��w��m�tZ����}.�zr�UTg�	]־pi'y�1hh��W)��궨j�,|55.�[��EP˚��Ώy��$��R�B��=?��� V���"[��䗸�hI~c��X�ny=+I�'���S��{�Gǽ]ϒM/���N�;��-�=����O���X���n���U`��;�yh-&f��MpIP�V�;��Q�)ۥ|!�p2Pű�.4�k�����)�I&��ܟ�$UV��9��䧮�"u~������{�o�u��%��`Q�_	� �Z>�Ew�*�����E#�r���lp>U�_���	�~,���)� \�-�RV��T�{q!��ϊ���􋠃H���������cm�ڒo%贃V�¸��&�7l��0�K��jK���ߵ�.G5|I.=�W�.�#W�  z|a�Ih���g�4ȋ����ę#�oT����[�~	w
b�LOUg{�-�..�������r9<o�߁~�X�����q]��s�����d��/�t��W{�"��L�I�2q)�N���r��������h�iQ��w���ꇛeJL2���IDq"V���M�b���9��ۏ���dG!�1�1���'qrk��A�¡�m�m\=HBt�l}k{_0G0���G�~�eK��q�a!�R{Z�h��Վ���Q:��$��a��h�a�?�ۜϘ�p��_���4[N+�=Oc7��0�h�z�)�$� ��|�[��	�s�\L�����t�7�WByx5����P2�hpJ����	o�E����迿A"�z>�� R��*�_�a�Ws�FCY�������~�Ԛ�z-�OD�b�;I�\��l��c�j�* �7h��2���������$��I���~.��CX�Rɪ+��,W�Sj�����pD&�-H�Y���F�J���)Wh��T�&��ڟ�Z�R�"�d0���:�$B��Wg�� �|�</�#]�(���� �ϓ�H�@��<�^M-�&7�I9J�3��VAX�㣾�>�����3���v�	��yC���f�;��}�g�a�ND��I��a��(�'�z��uB,,W����7���Χ�H7�r�}�zϸ��T=��(Dw��Z���:��Њ"
l� �����5�g�P����JBr��T_뷆w�@CxԆ�t�5gl��8���L~����u1�	�ጄ7^�AKݝ~Y�ڇkf��p�"�D*��2�Y܋3-��#j����,V�ޠ̼�������q�K�L���|�a���%M�f�:��g�M7��B�gsi���aQ�U�Q���(m�/�?е͠{M9i+S�<0�wW����J@]t�&���<�o�e��s�����p�H�+tp�����\�io��
�r��-�t��Z��]f�1��g�b�eL��K�W�X��0\��U>�� ��Z�ϽCR�ܲˣ�-�bMt�_pL�G
=�C���� zZnp؉���⨦'KTK�в ]Ic{**k%��F���y��+�(�|[������/PG��PS�K�	DΕ����^��<[�6��;i�6����I�����#��GC��v��󏖖t�+���%�PyF����ctjKu�+<ʖ���Q�N��c�gِ��u��(6�.����!���A!�Ί+���oR��:}r�����#td�Q���/_գ�]n��X	k&� �z�5Y�m�oRFR}�w��P�����.�N���fx"6���*�uE:���0�ne�=�Ɇ�e�`�x�<ӽ���/}�'��ɩ=�v��s
�2Rݲ�5#w3̑ �:1�6�U�#�o�	2�.�B#s[�]O�j�mh�dl���}	)c��Ml�K�?m����rb։�{� �4XT��̡{�TH�� ��#A)'����V�s�^mC���V�&?��r	�-�.<BiוDK;�Ӽ�%�<V芍W��9�*T��]7(��
GE�gu���2��)�	�R��7/�K��S׀�qs�g!�L�N0)����Am���ɖs?2���Yd��6������뤢��'�A\�H�[�J��ut��a�?��x&��V�����/�86�f!�i ���jG�烈?�0�Κ漚\��kreNY9��F��w@i� �x�xN��1�o$�@���ӿ��YU{��+B���g h��~�D"G}P\Kv}��::�*�ۜ�>�KN�?��A�h�Y��vK�N�t���7J�-�����q]%����ռ�*��)h�<��1�B����0�[��N]�û�Ra�%�O���cq`�(6���v��xq�����R�R�W��K������ڴr ��i9�'�E0Qo�O��<��[�4�=v$���j�X�ٙ�Ur[����'���e��s:�(��t�N֩7�\�Kd�`Y�5f���ZI� �f͏�������r������ v�8����t6��vY�qk�׈�����Z`��I��m�h�����u��� +���|���_��Z#���T�V�[�эyE�L3�i'1��f�~�z/�t��*����JaԜD)L#��[��9�V
i����
�B�|�]h�R����F����2�W� 9,��G�Vo����t��e�l�^����
/�>����`X��IX��s�	,��o!�ɱ�WV�:�KŚ���b«_�����_u�E����g����HHc+���-��y�ژ߸S��P!҇�	�IE��M�|	�s���
�SAgH��cZ�R�u���e�~s��Dd?"��a4^���#�w�$��tLd9������K}��;Iiރ!����c�Tߐ!��QH�|�0�u�L��������`%��f�럢m�3R�$SZSz�?^2E�dLX�_�u|�?wCrW'�!����ć!��u{-�i�|��Vm|�ȯs_��)�����suF���Y�_Cd�(�d�큰�򣽭5=�f�Zm���x�#*�q��C�$R��"i�J������ :��"X�"���{�M�-࿼�&V���<���jDG�/�v��Å���!�zQ�ˁ>c���?)����ߙc��Q�?�����1>�Fh�s�6�4cBX�������=�����L*QuȈ��Ƀ� >�KX���`�9�7������)���q��GďVLf:»m>�1Y����C_��z�|�l��;92X���R�r~����{ �	�k6�i�D:�h�u��z�:���V��e��D�ˮ��1��oXr(�#�υ���AїZh�9��ju.ݵyJl®C"�!��!�ґC:�VA��AM��i��'��C����DvG��C�]9)n�F��*�m��h�wRB�u�o3{h5}&�����U������E���u�ڄz�1޸{���@NZu�-|, GA~�%e���c��?������{d ��Q����%$�;�g���[D|��*�{=HQ?��'���
�(�/��Ž1ͷhݕD�}U����+�\֩RxdT��ǰ������E �i���΢2@Wx�YY=T�v�-�~��ol�/�&K���O�+����B�ׂ��O�bK:��j��:¶���C,�lU/�:p�d��ay���J�I6`����q�[L�K�tgo�<��ה�w��|��,?y�B�Ϡ�[��2��n�>q��=G�x�*�2��z��&�\�� ��@I�+�J�%q=mn�૷tfk5���[)F��LS�$0�	kaOl~�<���ԼJ�2�_��m��H����e{���y|hw͙9u۬�m�[��5�-��Ͳ9�\.��)�
��X�ݯ��Y�������z�yx���o����Q�&������;u��z�t���D�3�:2`(��u&�n���6t4
�:�	B�\;���S`G3`;��o�h����=2��CP�ܝ�X�7�
�%ؿU����f�lØ׈��7��M����贬 ���T����ؑ>á:�5,��Zz�Rݲ4D����>Ó�|N��Y�������;���8�m��gr�j4�-�_zܠ�(x���@�������U�А��w!�L�`��!�h��~r��^S�������qFP�)m%ˉU6��IZ	hq`����d�a��y��=�� |�4 ��t���g���g�+P&�j\�|2��멿�z�U�G��ˡ�>��)�-C�����OT�kZX�ɁH\���p�b
���0��r����b�?� ���LiV��E�L���!9������4�L�R��U0��w��x)p PC��ͩ?H���H����%����TjC��N,�m"�w�s�V�b +A�/u��� [�Y��������$�f+�\��&b�{��|�.�@0������s2ξ��p,5L"7�M�~}q#�3i�S���<�����/"-�8��ϟ�:�U<N��Q�d퀱�l�)�AL��ul���B	R���#����Ѝ/����}\�}y�=p܏K<'4��v�#�Ӹ��z�2M��H��ȼ��%?�$^c�X�'7�gH�Y�rjK竆ta���E�
�^޾\�|y��H�Xt�fK�ɋ���kG	���Bj��v)U���1�T��ER��_A(��+��3�l��u-;���44�h�h��� ~ �U3�iE�k���E�bm$C.K�9�d��ߗ$��X�5�_��_�"���� f+p �Bh2n��֒r�r��`���谭���ŝ�<�tq ������n�z�'�S,��R�$�v������B~��ٷ=�Sz�|��N�#����#v�$IBj�#�[W����[����9Oq��.�#��CN�3Zz�0e��SF��v�l����,�TB��n�(��5_4�eP��:�UKB*w��8�>��^�d s�e�)�s,Ls��\0xѬZ���� D�ܹ���k�>2p���	@o��'L����e5��)���X���f��6~OÆ�2��l=f���A0�$������&p�f��vj}�P1��wx���d���gv,�˷x�c�	7���'{M�J�+�r�?�If��F;*,d߳�̈́Z�?����J@5�э�Q�����f]$N��u�`�iv�Io�9�h��06�u����(R,WP/b�֗��"Ε�2��e?b5�6����e�P^&2z�& ���;�*"?HQ����HG�?���7��T��be���@Q��T5��U�߹ ζ�J)�V�OP{��)�I^M��	s>d�����o�y���W/<����ff9K�����X���*��#�O��!�#�N	�>;�*�Mt=��o���מ�p���tX�0��C��࣫�v5oNI|#P�A�6��Q��c�c;A�$���R��/=�^r��V(�;Ğ
�����*�5Bφ��/V ���B�5�.�`�#Ό �h$�Fu���m�:��q���e�0K;���z����ܿb �,��&�ǿ��.9��;Iy,4�A~X�ox۔��7���F�C
V��{M��w��u��V}8�2���������l��%!�i�`SIq�Yϕ"�'�)���J�#a� ��b��������qޡ_�[�6�ع\�p�ѽ��!m����P�^�Y��ɂ�F��IP�$Y��D:)��*�	dǺ�D�6#Oy0g�����Vo۹̏�"�b������2���;Ct���Ѥ�F�,n�u���7s;���t��W�8��~��E�d��c�@�x��x�Pt=#� 9�{�mp�2h	
d�� ;Lk2I���gW>V -�'�W5����E���f�2�\��HT@,H�LX�^���G=u5`~f��ÞWw��|���pl7�O���aY3��l��O)ʎ���BW��?��@������X7�×Vd�#�|�f`]�c��o(�s��?Xomm�� ������:"܆��.x]c�h�g� \��U�V��G��i�,�&��	5��6���~;���΅�ϼ@E���?\��{#��W��|��k�;��<�o��C��׍�h%��-$��s/2k|Vw������&���S=��y}x��ZXd~׉�a��p˄V8�E�e3����v��ʵ<..�Jov�R�H��J~�A�#é�A���{�)q�)�� ��#HS;���0-�3+�vah��u+�����J���P{���=I3�v����ri���/��=���W"��Ɵ{;g�T�`�e^�d�3N�Ȑ".�St��1L-�b�� z/�=;�=����-{��T@AjN~�
�}�o����gT�Ɯ�dи�Ur*������p����z���d3�Z�e�R���4k�,�D�Ɔ�78������y#�3�[n���Ō�+�%E��-j�W������+�r��~�,���t�:4���d������e�)�����ӥ�:�U�R��aB/܊��`��`�`x�xں�Y�jqGֺ�.Q�^��\�7�G���|����8�=VrPV�]���؏�UG�ٚ&��6q�~
���+\�]�(#�sBCpE�SOtuII�iʩ𵸮��t�_a���	y�P��:�u �RDb�HHxm S���JƉ���9���2EZ��Y/!>Z�C��$&�֥�����s4I�i0��F-֟/E���͕�p�2�G�4�^���p."��j2ƣ��� �Õu[l�K�"q[ҔJ3�0D�����s��ˮ��U��D��yX���9�[�U���e�C���1��~���BC��1z���ӄe��9� jￌ�ܲYa]	k����g�fDN�6����D��{�ڋ�lYѦx�d������d�B����6Pٹ j���|T�a����9�<�߸7���"�P�nP���}���6J>��A)6F�ZT6������,(����-�U@q@]�카���?�4�7T��Ԍ�'%I*�������z���T�OM8���k���WE�4�?I8�����]�K.S�V-)����woH����N��׭��L�5�k ����ϥtJƒ���6c�S�S�w_YF�ss	�^�6�Z�v �-�K7��Ǫ�N�Y[Y�*�BSwUE�X���L&,,UiH�fv��{p���3�Gp��xR��wz_L��D������ai�EF�� ��/sA}p.�i�a��P5�[&�am�,�Tcc
M�Q1#te�4�͹I�:ۊ˥.|�s�bZ��42	�[���k� ��$*.�o��������q��O����.eW���.<	�E�*~�'���T��
��-p�b�0ߣҤ�����)*����	"�6����_��d�\�Ή�3�^��8BW���2Dc��
g���KX��[˙_f��������bQ;lƖ6&��T�H0�ݳc oiOxS��v��KR˺���e�d�lM�APrUR�7Mϵ�)GI���s<3�ٯ�U\�foh�m�Ȇ<]��`7Vfq�H��
�^���w�h]g�g��Fr�,��W�Qv���st����a�ܩ��a�7���5r��b��k0�n(�#��P(��/�i��,HZ� /i>���'��u����zWP���O�|E!���jɈ��|�-���xva�E�ɹ��I��7e?����1 �I�Ȭ:Ux�Y@�lQ�J�Jy�̇3�8Ϙ��x�̲А�}��r^�E���*��~���u��\W�c�+��*��Z&F��[H�:�z%I���I�dQ�w��#�_��4�i~��:�SM�	&>h"�8BĿ\�<�wr�݆
���֓�L	�� ������b�n�Ay��Ϗ@�i���^ ��H�����!D��#W2�K�׹	� 2�o�A��@LT��=	�7��4��˚N�vQA�Lu��9����e3֌ �m~ 7�3������	�:Ɲ؂�錖�ǲV̎��`T�2Ak�ò�����ʭ}��9Ƥg>�L�kf�s�тa�����,;����<i?֔�/`��h�V�����U�YwuH�P��6�񓫛�ݔC~�O��Q�aO�nsQ�T"�@��6��w5`d�"e�e��61X�/�z*���Np�=Nϳ�Z}���̒�Am@�%��T�j!X��.�4�~��C~B`j)t���|�\��l����*1+��a]]�0�\ɂ���P���i�CK�r���#��p��\��Z�NJ���^F��rG� ��q�˃���H���=�����N%l�ꢀ2�}3�p�"���V��(�X�N$큰aC�;�]^[a��(�$�v,ښ|'6�Fve{qʔ�#׎��-Y�P��(��x�S�lѺ�>�0�{=�G��'8%����`����	�_SX?n��l"�__JB���_��_pz\����2Q}C[J�O���U�?���	�{��gYQv}�N�i�Ą<�u�4�?׳w8����)�;`e�T�s�Qi�~�Ϛ9�$"�#�r�R8�E�v�2��U��W�"�6�&
�u۵e%'�A��r'��h�A����˪7Cߡ��������4]Y-��u���8�^/�(�
�� �(�/��#Ҡ-��*(J-�t ��N�V'ȯ��+Z�üV�F As��ۘ�7�h�?eY�W�V�}GN���y��~@�P�.g����Q z׵�\GP�t���+�Rw񂗭RwYI�Ʉ�X&ϲ]z���3��r�rby�/#�Fy'30i?*Ҏ��J���V�8w0��˖ԫ[�o�ST�3�t�g�sճ��uDFU/��֘ݾ"��+d�Q$��nlF�g^�e�V�w�ܶ�1\"V����<�p�s!�q f���S��yKh��ZǮ�9f���qT�j&Tu7@�e:g��6��A�C��lg�2�X`-	���9�����!�C�춢<�0^ǫZ$�B4d̒r��6�����w�}�8#�kY؃3/�YINBj&�Ҡ�"��3x�G�P[hj�'2����q��Rt���292U
��-��9����Z�X�O�^K��+���I�G�����t����4�_�u�{��TA�E[��O:��hw9o�ӛ����J��1YK|U���yc���8�*��^��P�󬥉�x�}�}Z�"�k ���Q���-�&/as�K�7���Xkz��Ԛa���w�!�w��I�{�2�X��x'l���I�8K��E��?��	��L���cRK�]C�;�N��Wx�9�Yay����#�mi�y�#0���v`:�ú,%�+].qK@uކ �������S�{��6eKya�shG/�XZ-�����3�z?� .+h-.�C���	zq>"VG�D��̊�E�qvh�C�{Z����^��I������/�t���m��E��,(zqU�7�G��WM:#ъ��ek���j�'�r�ܴ9��Ƞ��YEN��{ˌ�SJ��c\d��Z�q� �t)���Y�s��dAh���1��Ҋk�z!�$���d���ە��!�JZ�+H�+C ���Xw��H8�Y�m#QO�)�\�\Y��~�ă�a��E��8��;rOKTia�4�����t�z?@��������s2�5R"YAW�:l���3m?�ﲠ����i�s�`�����Ob-�g���!�)"�G@Mp�*��c;�N˄�,�<f�s�����#˺$h��;W�ub���Zu����
���d  ���^�p���Kٍ� EMׯϩ�O���x��{������ ���̓���]S�}���Y�o6��VpEK섌���ia���\��>��n�M�W�ڝ1�J��Qݬ5����OHf �C>>�J6���S_���#k#�oC���e/��;��ȧl��߱����j�����-��ܫ�r0!wɢ�C,�����;w�8苆�q�#��ѱ����DB^�?�sl�,��T���8��H?RK ��e��'M y��ro�i�I0���4�����Y!�_�V!��n{�n?|P�:fm�#`�B�Q&���+��~߱i�я�3�kG� ���x6Q�0����q��A�¥̶2iW<>Rt�v����)0J�����^G�Z)��YdO7�k�����>���u过ڃ�
�]���>^�.��k`�tM�7�l�[ر�v>�@Zpapd��Is��``�o�.)�һ=���9��4	��z���,4uF�<ھ�k��ɝ�G_�
r�i��?e�]�n	R��2����\ցr	��*�.�/R�����.�?��B#%�l�����"����7�u;��X�5
�	�$D{�Z�����p��`��w�#o��o*�,-�]��f��ٯW�n߈�L�!���*�bY�C�y4�7�:�3$>��Y�"<�lE�+�[�wj����h�0R����L��W\���rI�U��+���t�Wem��D�7�>m�es�8i{И��80 ӗ\��e�h�#+�/e4[�L��FO���^��PW�-�{�Q��NR��Нw��<��9m�p����	���/�CJm�h:3{���kK�M�lz�izDs���&����j����Yad��}���&rn�_e�;A@�I/�*��m
c��<2�����Ā��/T���#���*�����f򣎺����fj�&f�ۖ^o����G�)��	\M��Ȣ'��7�Ǫ��P�� �@U��X���ε�.܂��ǈ�b���y�B䆹��8� 6��®�0M�k�b杨����s�g�4��qFxLF������Q��/�Fp [���"���k��YKs}�n2��`�89j�1VU����q|"A�D#���폋�o�4�1�9��G��Wp��@<�_6{�°e�ɱה�fY�,~��F����S�g2���?C�Tk����5�J�,嬍����ڑ9G��X���U�s1 8O�Xa���#���ٶZ�_ZUH��P�7O�|ɱ� l`�it��e���&�6g��Ž��[�)�/YEC�p�dh�\��N�|�x�%�}�$��R:9� ʷ��֡�KN��%8�1�||��Y���M���k��*G̙Q)ދy����o���kiQ��j�骅���/!]Zzj`1M4��@�f/r����I�~��f�������)o*ݶR��O�?K����q{��ԬК��<z�iݯw�ض�z��r#Պઽ��F�H� �Ş��_^$���훓���U�E��5��8�����A�k�B�� �3u���sV��	(b >~��3R��ؾ��]���*�ߔR,�����w�(���1Ī�z���9�A���i��KNC�0kI2`��?'�C��5����\�15�T	8�W#6���z�&��������$�zWb�}��V�I��N��
���VS�ƿ��[�˴�Ĳ�ބ&O8U��`�?�7VޚW����O&����>��'H_	��"�������z�=��j�5:�!�Z,<1�Gq�Y+l��fYx*iZ#f0�3�9 x���_=�5�T�*q�� ��r݌�E��cxoq��F�z�(�x��IF��GV��`�����B�h �Q�?I���Yγ.#�\�L�gy!f����,����J�����e�/N�ת!lT�>Y�$v�mz���P��!Sg )�%5Q��ɬˇ+�@�c�G���'I���M�e�03��mM:6hkne�D�������#4`�ݩ$m��j��+�
�w9�e�ԟ�.�}�xUJu�i6�`��	L�(�"aLS̗��"�w0}+0����E�����h��Y� ����u�msAȃNfkz�ɕ��v�A�����a�%�ٌr]6^�S���7+��~;�-��\���N����H6��~��W(C�4��Σ-��X����(=���vH�S�5Q!�bAinThP��F2xA�U1�#/�񄲘1�d�A�az�=���Ђ%^�1��׬�r� ���F��`�����.���#j��
��L�Z.�b1��6�Td��«^� i� ��#X?���"�<Pm�-���'U��Z��c>~��������cu9���G��k��l�d��H��g �'P�-�\�t�6L���Y�r��:]܄�óh/õ�����\z���Wz�a����H MZs�x�c�F�(gV$�f1r?��*!�X1J���ZV�A:إX�'����/I�ܒ�ުXB��}����
��.����P�$�w�4���� 4[��V/Q�z��;���Wg��ǖ[Y�����hE��π/��.ɛ��Gi�"��jVd��� a�����t��=YǞԩ(t������N��)B"��b�)��`3�夤�Z%q��`P,��ŕ{cj0����۬k�/r��aej���~�p���⍹���2����nYỜ��x"	5u�8���$nyVۂٮvG~��<sK �j�*�fZ��*ZuД�u!c+a�+8Vo]���}G;+F$����ɹ3jߏ����y���5 �Sγd�ř����ˎ�P��^~V�(O�G}��Ꞃ��~������5�(G�9$����*��=ܐ��H!�z����f������ž�M�T��{G�-ඩ��lj�q� ϰX�LVՐ%{�5_ X�	a-��3��㦗a�Ѯ����5��%ns��:r����Y&�v�I����1��_�Q�\����Mu������ħ���) � y����k#Li6�e͙�9&�)�Φͭ�����,���zl��V�n��6���W9��2��e1h�7"�#��Ɔ0���V�I&��{.f����՛�W?jV|YX�[�S�O��dJ�WZ��I������Ӻ([E�1���Ɂcv7���/��G�́^�����u!���]0F5��#8�_רp����5N�}��8b)耪�'E~��ӯJg���[M����kHb��3n�~U�GH��S��$��f���n(p �hs\��t��]�{��`�y门F�@QpSV�5	�[L�{��?����v����1�\<��Y�M�l� 
�a��#`"Od �z�D���q����㞡�.E
�<�*���~x���Jy�s� z��gh9R��7�&ӛ��WL�����%y���4����m�S�K`�({$>}鼔D1Ĕ�,nxs�/���6e�s��x�b���GX�kƠ�[ظ�,�����ũ6�z�c�JW�`���o�� �n��+�U��O�jb>��h���)\�r��x(En:�`Cq*_��L��C��e��Q��y�n���*T�%�@��C��O����c��h��p����z�]�7Ԉ�Y�7gݣ��Dڟ��G_ޘ��Q@�&�_@�6N���t�~����NSEk4m�մ�����	�z�!���H��j�-,	 d�0�(��h��r��Fr�k�Hk����&���U��mn�՝�@3����S
���ԿH*�	������cx�rR�'��[6�mG�a#O�ߠ�7�lam#��c�Z�~d�L=�i[j�8ug�ī^�]1�|���e��APX�a�M�,z�u���3�_߱)��$b�]2\e�+��
_e���9{����J�Q=�cF2j.�w3#��a��5y`F��>������P{�`�g����`r`9�e<�>)9G��k���q��|�+Rv�و�Z��KꪼcN��eU���+oK�6��N"#�`r�!��f^�葫^����j�@��r{�!qT@ K�)pp�*���!���E�[�>Cp�hڮ;Upk4�WE������2Ro�hq�%I��Vc"�_N�����$}$�_��j/>���1	H���C��?�YƠ�oW�ۧ�6Lc����\���k7��:y
8\҂�W�N���ٴ��m�tܺ&���#A�&�ALsh	U�e�b�K�N=���R~��m����f�$Gm/�0mIa�sG�D�b2�K(3�����]0��u:��q�hPٴuS����;�����
[�j^��P���#�|��ߚV��ڏ�-:<�3b%gI_�ۍ�Mӡ�ν7rA��f9�FD1�����S��Q|�-���0�~_8mzo,���&��Q5؎Z޴�R3�[`�:��1��A�%�o+6��U��̝�;���NI�{-�DG�I�p�ChT��E��g`�k��y����U?�S�{n҂�;��-d����n<��\�6��[ �F(@����M�j5�{ ��Ï�Qr�xD/�'旡�$t��|)W7��!�q���釺TJ�cсԧ�8cI޿U1�B���M7 ND�R(���_��ݐ��9	���[ܓ-ǚ��i<�}�9�I��Ĵ%ڇ��Ia��C���NJR�(D^K5,
��Z��{8��?��*;s۵�B~��L����L�E?9a?�0$���������~�'������?��$E}A{^7����O>�&�-���j4��#ӫg�y�G`�)�{S2R]{1#��-|f�����࿢���zzrU�{�}�é�;�J�ϫ�b�x���6yLE����K������c�|���~�D�\���̅ZD�$=���;3s&���S�W�U�6[-���aX$��wݳ0oҹ�L����qU�z�%��H����xk0e���E��@��)2C����lL�li��ǡ�{Ez��bz���כ�ө�>�lL,�~�ߺ�
��/��%�MG<�l�����2�D`	>�W;�ۨ�ť�4a( �%[��V��|`���d
R��$>����8���n������i���u'�_fzn�mW$Χ�1�uP~�t�8��\x��� Ud
ɒ�x�:6����]p�;��݊JSެ����h�"��L�7�b⠄zL��k��r��b_SX�%�\���eU��D��1�{�E�� �RB}j�ؼG�R%��Q���(*R�ƣ�j�vD�fq����=���K��5_i�UOH*�h&�:+_O��HW��y "V�h��C�F�Q׋Y��73�I��b�	���
 ���M�jqI�����CGr����G���$�C�Wʈ�~�즏Y��g> �Q
W}�B}�,��#k1
��n�a�੦�	�E����X*!˄c���lk>�{��c7غ_⍏Si~�G��=O6���?Y6ɜ��x~�Ni���gcf�� �Wǽ�Az���jƊĨ�,��E���lK�:���W$�Nr�`P�-^�-�Q�³��N��>\RF�#cLA:^?<��2w�On���a��9m�/!�'q��o��̆]����+�,{���N���:.����KՀe���R�Q�j���'^� m���\����`4N������X:��}����t�ZXX���H��zHi� ���d�����(���nt֝���"iDH��,x7I��O���`q8��k'��xJ|>���#\��V�V�gJ-�	9d���4_���_=(arF��[��m��n��M�`��r��2I�VM>����S��o�����ہ�PS���g�3�8�R��t�zQ/@3A�|Dt���Y�ӽsd]�����1Uf�'���0Rj�\���!���XoN��y��Rq� �Z8�>�A��z����r�\�b9s�:��G\�G�m��0�Uch����|\��' _�Ҍ�$�����+y3�֯]��4���ʐ�]is���W�>��s9�𩞷�ɄhV�ؒ�=$���W�'Ќ�eG<2��G=�ǂD.$��OJ�o9�c�i�ДX��Y��T�-������%0`��a�g�c��Y���V�5��3R|��gD���
��
Qvo6����/���lY��#-�	�PL��A��#��tU/�z�ϫ>�M:O��"q)�������}%ܘ�S𤭰6]���(7�:�[L
��hqH�;ӷ��x�r+')%z¶�pG�y��Zi�+h����l푐��?�h���GGG� ���QG��ͱ��/���$��iL������zh�M�4}�B��[l�,3�R�H&�O:�G�<Pȥ�bsJ���^�2^���?��6�,v�'r<O�ׅ|A�F<'����aV<%}��/�Y�����!G���RzW���=b����|����pF:F���iQ�izK.$�"Ͱ J��o�/�Z�u,�B�#�}!����h�e��%��Y� B������C�=	~X�z�9�ه,	�*�?��G������䣁��E��Q>�0]�y/�+p�-����Ѳ����2�mc:��ғC���X�����,z�կi���ְ�B�uh*�P�}��(1�0x|�~��/j�T���ѻ���\�$&<<�6v�������	�%��!�gV����"�2s��}��}7�9�*���V�cPr���]￺�6h�G�Oݔ�����#��x�|�s��ݤ�V�B���$�m����З|��<k�mm������A\I�f�/*�nЛ��IYH!��:d�ql�l|��Uu��f���>�w!'�`-��S�*�it�:���*F�
�����!6Đ&T�L�bQ�u��p�B'7�EL�&��|���am#�{t���j�X���F3\��.J�4�:অO�ܙ�8���"�vC��/b/�3Ɯ��P�j��i��d}�:=�T�,޴�dF82gh��D��i�L�t%2W�Y�T�:��]
4sY�$$�`[MΈkZ�M�Z%h�51+Y�$-Q�P �g\��*�����/!�A��8�@)�Q�,��⺵?A��h�͊��=�5ڸ���럱�(@���6�;�Cb�%^��]p���hm�� <��E;n�?������/U�*M�=�1�}�鵺,@u{��Lc<�	�_j|���ͼ����9|�䲨��K۠h	e&i�<�X���YX��.�����C �N��c�t��,$S�5�NxJ��W��H����s7��[���CO��?�x�Fy��)�󂯘�����r�tVb����5�Ӏ�!��E=��S�r�']7}�
MS��b6l�bp��%s4�+�lr�.�|�=@�ʤK���$zJF(���z�L��!���2����/1]��r�\$uN��h���������Tw�
�?�e���^�k��NHm���@,%=�s�l�t%���uu`��۱7��F�
���$)�\rz]O�L*Ǫ�]i��A%�%vi�)��w]��y���{S΋����O�����f�Ӟ�u�������o�͖�q㿰���}a�� M��D�	��tUm&4���!�;f�\���Ϲj,{J=�_�����n]�.m���Ar�j�@��uC�	E/k[�����i4� _���a�"&}՚5]��h*�F��g�ވ	#��k����W>��N��}�>'#�JӼ�;3_�W{u�̲Dd��0c�8�H���_���
P����ؽA��t2��Č�u�7)U�Y|m���Z���S�{~-$�'Sw�C�hui��fv�)`��~Gl�0yh���$�J8㓕��'�����H�u��0�i'��9|:�UWwE?j'R����9�_U��KY���f��Ȯ�xS@����/��e k��'��Pp.e��$�_���z�W��O�\���b(A�Nb�N7��H�I�EW��� ����E������aK�(���φ���K�����@ߴ �V�W�|�?x�έ��'l��o���<�֦Qm���>#+�ÿܵ��|�?��#��\pȫO�,���,�L�N�OMG�<�^gn@hݮ���{���pB�R�H�U4 \\��0��B�����b�E�.(Z���]�� Q�G�����U�e�-�����9�gL�w#�cl�~`�h�]����Zg�K�f ��K�.ջ1>2=�A�1�֑��CmS�ɫ��t.�0I�7ws"��I�<L�o̿��-Oc�֧/�$�������=Uz�#O���0B'�Σ[[�)����va� �~�|�+�0VǶp�%Ę�%��ք�5�˩=Ʒ*�y�.Ǐ�,$�1'�C.^D����!4�?�ް5�!�u2�ۂMv&��܇IVQ�տL~���`F�o@K��GB�B �_�ۧ|���ȟg
�t��#�>�獥Ps���R	�)�C�l�bSPQ�\n�I�Jv1��>��ʈ8p�)(ows��g�խ�l�E�>]�X��V��e���׼?�I���������7e�K�6��.�.�Q ����}�ά���J����=I��1��ɮ�a)��=剻j��+�T�W��@�f\A����^��2���|�9)�Q@X������3Z3�|����÷�����ƶ��Z�!J<�p�@��Y�3DS�߻6 }��9�"�W�E�&��䵩��bO򅤆Ap=�ٷ~�L)(vAܻK�1���j��fz�����PG�f���4�{/�;�V�s!�U
�º#
�����M0ns���P�VU�|�D�-�&��7߈���y���2�DQ��x_Y�k�%���*Y��(��or&*�Nn��l�v�/�/�2qH?�P�Ba��#�Cgy2���(ӜU_`�]�>7^
���V�\�9fO�+�|�.¬Ϙ\�ug����¥��z9�P����E�c��$�Y��6�544�lT�a
�,O!��6S�0��퉶��Zb)n{�$L��y�?M�E��"/vm�o�����������أ ��[~�F���>�*	�N����|u�pĶ5�r�>ث��mX=��9�����E���W�����@!)�oOj��bL'RCT &�h�����A����&7��LK���&a�3S�x�		^��A�,�V:�E��V�R ᤬(�fy���;���O�g}��n���Qw�ĳ��h�e���?g+���k�Cgy!�ΠX/\9!]h/"6�j�P���p7�q���j�L%�.�b2ά����3�?µ�ҩq7���LU3�kWLX��W�
^t�Cf�ߣ5��n��p����!��>(���Ga����������zW��X�!�|t;}^"X|*��95ߌ������*CpA�A<�GC��P�R� ���߿�"��$x����m���3���ֹ���%B�/ kv���8и�C�7���"�}�B�ҍ���Q�_�>�1�-�-Ұ{usZ�cY!L��M�AA1s��g/��D�g���h̞������B������K���e�ͮ��50&*�֜�:%��3ie��Ҁ�����B��P��a�zF�s3��=��T������mk�X��/�5�Ul��z��!ݚ���%&���-���ً�Oo1	���Z.�a-݌��B����������VT�uֺ�v��F�s�7D�F	�Iw�^-E\/FMw��"���bT��{k��F|�el.D�]�=D:�j��{�!e�A�Yb����@�k�M�\deï�
����V+9,+̶�d�X���<��\��d�NTh��L�'(�`\�oz�(}�ȅ���������
�;���vP���;�K�!|�+���Nڣ�G����;��!�P[�Z�U،{�R������+���BWL�ȓ��n���$]?
rX�䟷^B�B#L�н�6nI�$&��+�l%�xPEO�5_�yú���vN���'y�>�+	f[E_޳k�8i�Ծ��Y�Ai,��W@Io;�����* ��P����r�Z��s�m6V|�D=�v���V��*Y�d*�J�B�c�0�I3�ԓWm�H�̓�D���E���q����$qǛ�D��g̀I��'�ÛEN� O[�_g	ٔIAm�v���HmW]zHa� �g���4Wm[Q �;���2��1�	R��T	���Z���F���c0�R�$���������Ye؁��z>I���z�a$b�	o?���|� �w2��ݸ<4�C�.��E=�,����;�͹e����R[�
#���e�����.(xۖF#���A-��Z
�0m?	��nla4	���L�UGxNʥ���J:�#�d(��2�OXF4��f[c�OY��A21�K�~�@0_���XR~#���ԁf�E՟�x[��վ}��&�z�@�Ø|)ܡ�E�T|���#f�e�dt�
�&�n�4���?��J�_F��Н+�/fj~����� Tn.dh�%�R����kvC5�2��y�M0��reh��I�Š��[1.GH�1���b��tBn<��"PX���&|T$=��N���Ss�2'�<P+Ё�e�Nh��p'�;��s,��>��d-vk���ɕ0��P}V�3b�y[�1��I��.u�U��"��%T�f���u��B�n�7Q)V���VL���+"�[�p=B�Ĺ/v�_ak���sV���tt��:�	�g��V�I�����ƞTd@��i�VZ�H���𝭃?u�4U'�X��L��UO�7��w�G;��%��=�_�5⇷��ν�#���mg�^�aj'n!�g� ��<�)�u���S�e��,�?�^ڙ�
��W%�[�w=�$�^0F ��Y�Z���tjZ�J��W�õ�U_t0'}p/$F�3g�dN�ؤ�P�~?�!_;����ێ�_��]�ya��KʛA������mLJ�b� �����࿳ŏD�H�
��Zom�\�r�3��5��me1�>;Łj����j��1<���<�R�d�u͊Tiz���s"���(9Lu�P"$�dwe� ���6x�,��>;dB�.��[5�����:���^묹Mt,f)B</�x��WtՒ���K�F8�e��jT�����ō��-Q��3�+`��B�����2�Cr�K��HM	D�ǻ�M���ݢ;��jlm=J�RS��΃����Z�Eg��`�\�ŉ��Kɧ`#�Q���xWh���
�_Ճs��o���E^z�� 6y�G��;�dg��B�4�{	��㴮�W�{K2����j��(�aaõ{T�F��?/˒�;p��UߕMϮ��7r?KeP-�.��@&�Ҽg�Ƃ���5e��`g������N/�6�Ax��l��%x�N���� ���I��9���8m�E�6h�ܜ4N�@b�w��evx
|̐���^�a0��q��n�i���	���	�=�=_4Mf��|߃Hl�	��_'BPU��(i�U{��<rI\;���CM�-��ɵ$uA��fԾF*o�OIfx��"b���e�U��M.j��87K�n��;{��X�V��v!zJ�{#"G�0��ku-���-�Jt������y{9D��k�?/��k�4��2f��FG�ǒ�f(�	����k����Q�r%��B��B� ��ê"}��.�t�[W� �<���^ў��}�#a�AW6=S6�t1?�Z�Hc�Y)q��j�EP3X
4���MJZ�G	��z@pڷ�E��9�u�4Zvp�vR��H:Wj�+N,�#�O�]w��49w�<WEK�r�e�A��b��/�R8{�.Tdt��sӫ�e�.@(���BL8�0� ϝ�z�t	GB@���/z�ܿ	�b��D�[H'�Ynu�,sꊬ�RC�)(=iMQ>�QD�<���ʶ�m@���I/��G9��&�?3^�!�L�zjW0cy��j��&y>���;dV��&[ީ�ABi���1!	Wt\�d���(�9�KcT��uj�V��~O�ɬ�zrډa8*z��/��w��݃í �����@}�=d��ޟ6�ǖ�\$�%�/A�.Ւ�Xt� ?�ⱻ����T��J[C� ���n,KN��;%H>7t��v�M$�Nj�Ґ���ӧU*@0~T�?o4İq��<�r�����0>��Cx_N�z4FbF4q����|S�4�O�8��qK�yaɮCX3�пI�-Ծ���22���n~��i����{$.ُ�	�B�II����%���̾[p�/@�~����{GH�p ���\�������T_k���?`�. P�T�Q����I)�����.DF6� �_��g�D�2]�	ӏ�#e��Z�~��L" ��aa�&#O-��GgR�(�f�0j������ V��/Xd�f6��	fa^dN�\i/�����2+��L�իu��8�S����=n��Z"��!��%�a����n*o��ᕁ�,+�������׾|����8B	~��y���i�wX�w�^��'�&N,CY��.:�	�O�&��#N��+�J����҅.	�C1` K���@��������l���k�Y�{iNx�D
�k$�#�	#��ݽqJ���;&��YF�I�6�.��yC�;��%KWOp(JAT�#�-oM���l�޺�(3�ֶDR@��O3���B������:;늦�����:�#&����6�d-�l?p��9v�Gn�r2�0��=��	=o.*��~�q����6�
R�\V\�
ֹ�U6�]��?��@�w�[qj�ʛ7MU�ԋkm9�Ӱ�}�(�O"S6�/�Oyf��H۫S�Ɇ��GU���<0�T.e�B� �<x�=���h��9c"��"@D��0,l#v�8��=�
�����ó䬄��Ȝ.�r�;G:�3�-���N��t0s��o+��W���ʝ.�Kc��V�������?�R�X�2�@��#��-4��DA؎�e�^~���V�R��4��N���#���;�贪�����x���D�T�vI�hu���K��w��8�|�Wwz�8en���r
�)9����j��h$�f���������&�ͯ�K@iP]��	@��T&����4ģL/8� ���1_������qH�:������I���8��P�I��ǉp�<�G��j�+�V�kz4��p�0+��yG^�A1)A������@o_������>�V8Ҕ�!g�v�K%�O&ȠL�*��w�����Y3>=^@�::��xkV{���b-���J�O{�%x^LJ�}+ngK$(B�u�c�}Bn\���ej��ؒ�%XJ��iYMD��3��s1���s�+�Ȫ�Za֒y��p�,�F����T�FN&�y�c�|g��Z*���T#s���y��L:���.9���}7�66R�l���<G��uw��X�ڑ�,�\�#fҹ��(�:5�ɶ����P* ��Ip��V t�7=�9�D������0��C|����YK��Й��O�5͌����>�Ô���i�NC�c=X�F��I��Zr���Ah�\D�Ǐ0�|T3��5�`�
P�4���SMx�*@����	9��;�b
�Ksͣq_̮3�-c�iD�11����o�eLM�Qٱ8d��벇�̹�`�+\��6��]ک<l-��DKhR��9Kq/$�HG��vJ���e[ �)�`����+'������L�ZW���dx�)>�l=���t���P��Z`%��>P���g�u��*�GUY���a�Y\z*�ڜ��,_תY�>��V��@����5�n=���o6���z��Bs�%�<{c����'T��﬚�'����k��
n�`��~�|� ��<΀Ɩ\�<���ņІ��И$�Ec��r*��37v�\�V��G	�N۫��>��
s&'��T�>�ﰘ��ܩ���ں�ݓڥ��N�X��j�.��~�O���0P3oi94a���V���Q2amm���
䗞c�fE�Ԁ�D=��vx�VY�6^�Z�6�|��a��$s#W*nH:��t>f���J�5:�O��?�w����o�^�JL��,G�5�q%��)8v<�7�P��ßT:�1)w���Q��9	끛�_՛�8�"������p�PG����7ZK�������
N���0[%�y�+�P���H
TV���L���BF2��|����T���ԁ�+z���3N>�0��z��ӿ�\�Ļ�gD]�4�k�u�U=m�`Z�����������S��C 6"�x���*Ӈ`_�ǜ�D7d�Q\g���8�H�z�|�AVL�41Zm����t�@�6z���-�dX��]�!�%��1��ys��&-�<[m��a�k�W|覡���L6�jC���H5�p<�;��:�QM�wз�T�l���2�ǀh�;}`�7��x֒� fc�	m,�g����ߥx���נ
�@g�����������rSh~{�CT	o>n���|EL�vi)-����V�J�,(Q٠�4�V!kA�C'����	������2�՛��YŊ"%XЄ����1��A3�@��I`J<�k8.c9)y�v<�q�^��+U#$MS���uٝ*���`�|%*��iȧ!=^s��fu��[�-h�B\h����3����Q���9Y
��iJ>�n�5�뱅"�����h�AN=yg��G�;[�v��.`%ӿ��|����.�?1��~q����o�N	Ԇ�!���v��LMЂ|L��<f�B���F��p�oL�I{O@(y,����~p��E�-�X�c��H�	%��)�q��1��GH���D�G�$*ne�i�ъ���r�y���"�;'��.�v%�{'�c	�s��0���.T�,�M��J��.p*�76�r�sA*2������ v��ɒ4႖��m�!غ5\��8FTC@�GG�ߺ/�\�9���OD!���t��
�g`@�Q�A�.,Q��|��Cu8I�js}���Z��㡓�f�gUĒN�x��C$N��Y[��xH���,~�w�(ͻj�s����v â�R�I�W�����YwĞv֏������ۺԺ�m��GK8�� ��m�=���Ʀ8x�8%�r���q�[7�� ��%	;�W7�qE�f�n��(1� ���8�%
��v�����Ǐ_���Fj��J��eD���8��`�mhMd�\U�eA�4z��>��pHa�j��%1�>�0Z(���25a�r�6|�:,�ZM#��NQqˠ��㎋�Ģ�4�g�f��*�`I��E#�k!۰ki ƄZ�G��߶�c���v�݊WX7���6j�0�f���)}H�(L��Ǥ	�V�8fq��>%���=5��I�y�y��Q�����1y]��
Y���j[���d�@5��2�Z?�hY؏P��M���'�����ү��|����^*�~�������D`+�b6ζzUA�T=�N�Z�*�#Up��ӑ-��4_��	�O�I�x�g���4U[z�'\U�q����I�,9�Y�Lb�Wy8q�������'|����g�L(C��@X4��IQ����ޅ�j�݋�G�����,'���|�e-�1]=��Ӫ�����D���Ӹܬ5���
�*���"O[��AJ�1J�7=/-a���z趀�!�!���&�%�ݏ�"w��s@#NڈJ����U!�c�>����A��P'�˻U�:,�>7� u�ek����T�3��J?���%`r`��LzX g�{��Т��l+(P~���A�WS9�e�->t�Db�!�=�'^�����KRbʋ'i��CL�`W.�j�hRF4Uc1h��y2��6���r�E�Q���@l����{1�&�n���U?\��A��_^1��V��D�|������W�u�D��B+���	r�Fp����O�Q0�bU.�?�K9�ɭ�����8���%�ث�{�Cqw*��8P?jCAm��d{����,��/:���?��Ǔw�9��K��L�5z*B���,^�T��b��f�Ega�:� y��Z�u-lJ�p�{�x���v�ؒf!���j$[ˀy���媶���8W,�ų��Z̳�����ݴ���{� ��yxUd���a�WW_��1��p'�QG�բ�(ۻ����9u��/ث�$~��P.*��z ����j��QLP�	���#���dvj��惘�߼�����$y�3�<�	b�Zc��O[f[��6���)�c�s6���������᣶���seQgeVY@�/�����SB��k�1ݲ���?�u�l��I�oȁm%@2��J��Y"�c���~<#�ě���ˬ��Z��|�]K{�K<�	N��cZ9�8�1��GlylݴufK�K疀�[�j����b���@)�݋Y��J�eU�������3�o��g~�wn�*ϖ��s?h�a++�~)��r��*dDy$��c֛�G���|�7���V10TZ��{ '��*�#�v�_бU�����CR���	ۈk���EW�ҏ���"�}����r �Vʹ=Ҽ��ɱ�I����w]���He
���Cy4V��.� @x�q�Q�U��Tl�ՅFi�\��W��.Z�h|$�k�ZGvT���%��3����Xs�'����mD�r�M�i�iaҴ�Ư�f��ҷbʕA���='z����mG�p�,���A�M��j����Ũ�;��2�;mH=���4%�ڲ��
m��S��
[�7��wD�D9��s�MU���u#�2�(p�{����,�3��:�Km��6��t����W^$��	ؓ;!�C�m|��<�[یعT����o�����)D��GW�Q߫{���G4
}Kp��K)���u.��d����ɏF.c�{�>��h��ʱ��3g �+~w�> ���Nii�^�𬓶Llln�~}���N�E��S�E��,�`�/l�4���>O�t$U�£�r�ќ�PھQ?	8�iS5HюۛRT 1),��P��ٱ"M1q�Ʌt`�+����u'1]p=��>���o��dp�|*�f�27B�=��+�O[��m��/�R�m���c<Y�W�|=R �h�T������"OR����*Z�ڕ��q���z�<�'�K����z���Z����֎�D53�AV�=%(L�ЇZ���>$�s�I�i|������W����?�x����fJ��������m�94 ��Ovcs��)T�� /��+���&�oO���U�<��R(�c�s��I1�*"8��YxE?D��f��jAC�U�b�Ӈq:F�����\!��ѳn��oV�'-ے#�)���$م��M�A�r'�:��ʚ��5�� R�bc�ZI±�z��ɉA,�x��YE|+�f��,(���E��H�co|)V�z�E _NuL��Dks�<��0G�dJՕ��tW�* ��X|C�Ϛ���� :Vۆ�[�-_~m�n�ͨ��<LtD��X�y<�T7���=��z�����U,�|0�QmڠKgƘ���\�����f�
勂����0�C�Я�t��zT(��S�5?]���=�#p�_9��t`�T|rܾ-��5mXq#�����L� /-����^v6��n���*���g/�����j\��P1�D�J�L��]0i�@R�f�˻1��Fi�~m�g6B���˰Qv��̑%��x���Ӥ������Z��6b�nV�Hjd�V�q�����o%�%�Kc+c�z�vs��ǔgǦ��+e�c�.	�G��*�p#�����tX+�3��;�jcQ�����qR��0�:�Cĝ��D�92f�O����H��U����UA�V˃�B+2C�%DD��>���D^�����ɉ�(',^��rh����r�w'e~���#[U�Q=K�:̟z��',<H�O�M2ȟ���9JQX��r
B[��<��NK�5M�[+�S��� �&����J��>�?���ᥘ"�x"vc󶹓ܲ��.S�5�����h��b�+4��ٗ���RM�;s�ƸDIQ�Ng�а�W{m�>,��1>�	�7]��/Q��Z�v�L^i�= $V���7 �3>�`v��Cs`ɐ��E���c�t����4;=��!"��$g뢹/��`�����2�^I���n��� �ﵲ������ڥɋ�>��S�����x̒׮�peQQr�����^��'��MJG_�.ّqD�@�O�9խ���W[ǝ ���������Ϸ����/��@�XQ�8/���m�ZR���6_f���D�J���އR	�j��O��y��ʅ �����N��mr�tZ���i�5*�+�F�!U{��N0/%���u�G����"m���1�OWJ�8n�y�s8?o2+D��3��'0s
<Oi�bxg��*��v�΋�!��$IU�F;+:��ƶ���B������t�K(��{���dVC��y��;�;%�_��թ���vO�E��h�;`�WA:��(�
���ro��O��F�0���*��>��^Ԯ��k�Q�ކ/��}*D���ߌCպ0��Wl�����r�/Q�BX�)�I9���T{-�yR���Q��ɔ���CW�K#7 v�?�ɓU���+FIg_�@t��61����m�V'YL �@��=�r�8�30K��/+��s:���8 Oǜ��U�ZX}~�N_khϴn����.�/vX<j�2\v���'NJ0�3��&��wDe�0z����&�}��+�@�Qb(m�ڴ-z�{��׼f+HYDw)�z2-�)�h��<��w��$Mo��]�G.���[~af���Y�"�l��D�����Np|�����Hgyۙx�zUg�	u��N �J8��7	:g�g�B���S�2[L�^U+�<d���0���@gL�S@
<�z��'|
��Q����Ka�!�f�a���C*��[q%Q
5g�[�'0&j՝�	2P�QL�|��v��-����a�id�jP�;���U�� l:�x��H�m�LN�������yKڮ���Z=��yed�Tb�x.����Z���8y�"j/���Z�K��F���*���x��	��=}�b�+#\Gt�5�I��Pw�X g:;�W��_6#w��ی.�����aR+�>�����}�Jw�䴂 �qF�+��B}�ɛN|d�%h�֎#���i���n:A�B�@_�do~TgVq�Gh���,��ܺGa ���*�,O3r՞:T������D/ӭX��LWD���7��	=F�+S3Q���Q��aG�w��듡Q<$B|҇�5}���92�:���G$�O���)A�����'kT%�+$+0�:��2h�1����]�?B����c����-^s�;?�v���v2B�mEj U���k���ѻ7"��d�D7�jv�E*u��� �1�&�p�Ȋ�s�N�H�� ���9N�$c��5y
���9�0b�ϋ��v�m]��������,9i��)�P�ժ֫{�fAu��lKS�+M�~�)���g$�O�S�ƪt��W��/.Ώ�<m'أ+`���R�E�C���҅Ȝ�օ��+1d(���KUNA�(@v�4�݇%v`��ݔᗁ�=��I�˕�� M�?.q�ֳ���ؠ	���cQ/P�{c���e�:��_��c�UY�A��^�Zv\-� �h)���"�4y׮��)]��hcW��I��/�Ԅ"z�-�k��5!A��G����A���B�,O�l�~'|�zQ���y= �A�w����쟱K��p{��h�����`��U��.,l0���J��w)��T��+~�]^��#a��Ů9Z�0wh���+v�8;&���-�Y3���������OTz _DB�d9�V*Br+]������SҲ	vŝ1��F���e���<?��T HC��&�
^m�K�K'}s�MOb5/�K*���
I8<5��z���W%�T?�e�V�o��2�
��y&,����p�ऐ���m��
/��L<��i;
/��a��F�Tr�M�x3�a���T9^�.;�AZ����A��s�u�^�e�`lu���0���RV1��������~��]�����߉�az�.#��(e�=D� ��_�bR��/R�|��[!p���éGx��R�w',`
� 
j���gA,]X*no
b���V�b'�\���y���!rs��ҙ<K�������ͪE�s�h��ڽU>�i_f���Å�w�m����t��E	*,5[=Ei:�ܳs�`����!�q�%�9��ICG����ru����C�����am���,F᥷���R0�����I��aRO��ˬV�Y��=�P[����@MGH8b�H�#ˣV�J�A��a����x�b	M�ƃ^RT�}�3��A+k��ZCoǳ���m���hW}3�����aC��l��Q��r2�%�6�L�~z�>,�7CM�l�B�5��է	�f �&�B�5��@�����(M��@��Ex��fS�ڋr�K@I�$G�˼�����h{&ƣF�Dh���ϖ����k.����H)X�m�iI����kM�_���&�kXA�"�AE�X�r��D��q�`_o6[��[��� u�ڤ��lu�Ǜ��a!��tJ(�����p���E�:A2o�Ɨŏ���>���X�J1e��O�	�[K͍r����h�,��0�:�֮����G!��UǓ���6��(�YY)s��c�ÖO�_���k�d�c�-��:��ڟ����dŽ�BP��C�nɴ�[��RP�)6�
nߩ�F`���URP`�o�����@��ȩd��iI DQ)܋ih~1j�i������RR씭}��Q�Q�{ >��NZj���|ϼ9�t�-�T���^e��*MP�n}B�Iم���,��`7ٶB*���+��l~����V�8B��Hb �,9"��l ي�M��\��i5�T��J���UT ��R�{g%�&��㴆p|&j�X��_ VlEM�y��u���t�]+l�Q%�P�h8xCZ�K}�f��Rq�$8�X]
�*�?G����2�1Q��2�l�
�`C"&��Dˋ6c�ʣ���\QU&��Z-%��6����S���Xg���s��3w��P'ke0��@s�K%�����!B	�a��9V��Dc�w#����h��Z��gk79��쓕m�Z;)R�x>S����U�M���������kW?��m��)3@w�;*�IQ�Y��{z��{�9AOd/)�;6%�{�Hm,�Oq��"��-s̤t�9�����.{�	/������W@����o�Wi�L��a�Ev�kX%Ew��G�<���s�Y͎L���q���i�wu�^��p���M4?�4|�s�n��ڌ`��(�����,&���/1����_h��#��jr!l��h�[n�+��&!"8��=��O��=�H��`=8d}��V�Ss�j�VgJl�zl��2�Ҝ�����ǃ���8��T$Z�E�M�R����
?�F0�Q�®��D�v�[���.;�{��u��.��O�i���s5+*KU�.6��C� �,5#k%G��t�v�ޜ<x���2����l�5S��Zt�<%!jj��秹d�!�=�h��Nqo�)�%,�qo'�#m;2����c�<���r�b��u����T�[�ވƮC��tO�>Vn�Ie�,|TfR�vh�7��p ��;�2�������~"�-Z�y^�x|��K������B5MO�����>�'���5;�D���0���,��;��v�e��$e?�[�_7���\�Iu��(���9^��ؐ�!�88�5��M��lz%t����)�G�@=�N�7X!pV���<3���k,v���W��U,%3����yQ�������{YE`��Q�!����n�Vo�Jd�A\����Q���
C5#��=� :���8�鞐�cO�'&����q�.M _)�i�����D��� ��ڣ���ѫ_�2�tM�@�윒�;�:hSIy�ڄ6n���i���TD6�4W,�u�8Љ���_P@�3n���\��e󀣦@���'/��Asc���RVa&���4�(N�%}�jT��s楮�������%�ꂌ�D�X F�<����R�/�-�n�.�
;���ߓ��d����"��?n��]E���@>go//L�ə�hrJ����W�%_�8�~]颊�wP�?}��O�<z#:�Ƕ=B6� �R����5���i�w�n=~	�جo�\I�>'��d��i,R=�R���t�n�e4��G��@��ZW�4s�����i����G����Y� ���c,u������urP%���w������ZWU����ټ�3�tl�	d�� &~Wة���:�־� OSX���[�3�QW�b*���:@ؤ�W�iDt�9f�{���*��-�L(�Gf��[�-F�n���Zշ�M� �9)�#��s
8����7C��dS��B�q�q�q�<R��ռ�d�F��X�6}��O7Ca��Vj;yF�Ȥ��W�:�4��<��8!w�DSQj'�3�HD�R��gm]&Ȍ�}����_���L�l��F#r����Jr*C�=��O)!��t}���U�����#���9#��۽����Á�?Š��G ˇ���CT�4B�ެ�h(1k_=��5��A%����-���jO�g���"��p�I�S'a��2�JCK������ҁ�^f�,�x{A[e���.�X�*�$��*y���X�ջ����[z������&�� j���_�~L}�E�3�͉�O6
�3v�DB,i☧D��12P�^yt�f�6an�6z�|��7G�
�&�^�3��m�{=v����d����ˌN}�3�)��w���ٶS[XYa����>6!;��q����;븢�Š�8���L�bc����D���l��``3p�Չ�e�G��sQ��O\�l+J�� X}�&Y��Ly���P:�{�C�I��9�����	��Cm7P%�"�j�t�(��VnY68��֑޿2�JN4#�Dܺ^��N����|9�U�� ��Y��:�Bu�I�U6�Q�~�q���"��1����n��Ei�O���-9���ҕT^OoSf���5��8+"��>/��I3�)�V��()ヹ�r����䳭ז	C�K-�c'S�LX��g�*0-����.D,��Og�-���
ߥ�X< �&� V��ۥDq�C �ά�@�e��@'�R���R��E���5<��k��\�k�[�v��g{��aei'�����W�9Z�Fr��]����.���b:�+�?��a�d,�[��-p�ڷ�/�se�+Z�i�	^|����I�jP�j&�L����t�~�\�����Uu.���z�Xn�-u�9E�mA������ON@g[��������i�d�,�x��f�hZ!y%h�&0$��[��������oh�7���̑��-�y��岌��N)�Ь��OR�������4_�����Kګ�a�jQ,S~��<���4F�.��x���\A��4.~ΑÀ��ݗ���ჩ�}`C�gD"m.$ą9�1����~��<����`��pye͟(�l�;���Q���1J���mF@PC�HN ��"~�s��l�Z �|�!@+���騶�Z���u�A�3ƫ��E�o�������k�B�&�J��;akR�@+��=v|t8@�@1�I�H��,��cBj}�^�`�Yi;X��s�I�J���~F�Hmlh
��������yP� )����R�vbj��j �W:&�d @�����%��J��
�Et0��ǽ�:��ޏr)�Zh/�dr��k�@Q�]��l���U-��i�O|��2�=o��~hI^y���ׯ�Y�頲���^�-Z���K���d����I@����=�D ���w����f�B����#i#Gn�HY�C[�3ӆ�p������M�m'd���gM؅��}�*����i��"��㷋�_���T�O#�8(�c��*�5a��"nJ9-ڌ�W��{�4��_@8�e� ��~���O��E��.+�䃗_@&��)q��G���1�.��M��g��ƽQ�ݻ�`�����JFͭ��q>"our��f�I�d�M���S�-��Tc[����/�y�rڞLܝ������vz�-/��{I�.c��u����H��ȥ�#(�,`o� �[�����<�6��������m�����I¦�":����+v�4$H{�Ъ���vXHő�hW���;.5�HSw�j���U��>��I(D^7c�n��U%ee޻_�U3 ?�����U2����ݽ6KB��f'�!ٞ�L�-"�U?�`~oe���G�;�:�	�H/}�q��u���:��/	�H���?>u����.!f���M ��tQ�8.II���F�A��郬1�Y�M��=��T�/��`�	�:ր��cЙ&���YL�]������(�+!]�,��k�ɥ闀\���_��~ Rv:;n��iI�ĸݮGA �!Z��p`3�i:�ޚ�
�\�]���r���Cq5
d\@��}��9O�΋3��a�p�Z�^��D��LrlpZ��&�l'	�9a��.f"SD�v9�IDX5��=m����$��b�E0�"x�-%�w$I�ɐ Ү���\('�2&��s'9h��(6��b��@��j�;
S��W�bK���4� ek��ҷ$Z��!"�=�J�N����K�^х���Q�l�b�wMʶ�8 G挼��ݭǨV9�� -�a�i�!��3ٕ	��	k �3���H8�.��/(|9Qd�?
�:�XuJ�Li� ݶ|���黰,�S.l����Xj!V�o���;�o�ɖo�5�����F�ܘ<�c�A�,�󊆙0��3��6.���h��JH��ޒ�8�ᔃ7��HAX�S��|ecN�oh�̚�9sM��Y&J��7�ָ�#x�H�B�1����S(��Pl����$a�� \���]���\�W�D[Q����:�
.B���r̥�����6[Z�1�z�M�@{�>��a4�4�_��=��Ee��(5�ы�����%\)��r���^��3�T<*�ݡk��?u�����7%E-'d�[��0��|y�O��-��+���m6
�ѡ������`*Q|[i�
�/YNmR�����!��Q�W�K�Y���W�Չ����*��B�˔Nꂬ-;�3�xM�a�#5L��e�`��Jӭ��;;KwJ�F��)�M%�[�
z@e,�>����P�S�u��w�3l�v|mUDp�2����KN4M��㚏�ooBq���ƖA��٦�@W;oi��o���\_\�3O������%� �����*ҩG�&Q^ۢ�G�����o��00-fx�yo��5��5��՝u�������ב�+^f<�k�	>l����ͺ
�%����JJ���:�\���6�h���/�����yO�9_/K߲j��1�{��[ �����%���+�A�E�sP\¾���p��\�'�J��>�M���0�r�!�5@�BuK�Ч�O�T�CkId��)�Q��<� Tee��B�K���+e>G#U��c.~��8����9�?jg�8��sQI�S�a?Ms]�B�4�du+�S��r�R97��NYJe��)Q�.�C�`�����=�V���d5�뽐��3RQҔ'�a`icĜ�5�0@i۷0���)H�'�����0�B�St��x^��ǅ4y�����Lfg���7��������)!�6����ʸ�)鉣��f����G�K����	��� �(�19�D'��ϩ��Ͱ�w�70���x�o5*�{��E�[��#[��S�;5����q�ȓ� �����)p.2rv/�H�8d�n��[~�*�R�W��
~�<r�8FN������t[��-[6\V�C4����a�~џ�������.�h-S�fA�ɫ��˦���m��N���u$H2_{��!�+f{�9 ��O]Q:Aʸ��j�}�Ud��kTs�g��/��eF�U���nj�&�<ȓ����i��}���K�ron$�L�TR�V��Oayg�Q_�2���Nr�^"��~�zq]]��Q6N�s���$�o����E&�ˉh i���fN�.�!s����pX���^�
��0E���s�>� 3�������W����:�A	a����I��R<�m�4�hY�B�w5��p�Vx���]�]���2o�Zj5��4A�[/�P9/�𿪼^m��$�`��h �h�s˴O%�t���)ү����õ��h���!v>v���n�B��j��&��x6��K��#7�Z\sxx�Ύ���/�w6Z2���n��2l&����ךk�-�(iҾ`u4İO�"�Y��g*b�$�I�cm�����I�� �|����'�{抪��T����I����t�XS��N�K�E����Y#���i�Ƭ��g��z,b6�Ǿ]�⹰j�F��8��K�q���9z�5�ɟ	<�d%ˢu vv��� �roc~xb�*�e��AK͐�#�E��#��Á�Ɵ���8����o����mz8�\��E�7��Ez?j~�ǧ6�H��F>l�N/<����?�f�Io�U�ACN��Y	I ~	ާ���6��9S�EX�o�Of��0�d�B�:����&F�	���[ЫFC\�6�i�"�z�T =�U����F�h�
�����$z5Gv��})?ȇ��B(*9�^g�8w� ;�A*���J��ԃ������3�7��[_�!��9S:��s�6�B��:C��+��c��S�+$�[p�t�$��R�n���3��I��3��{�)���U���%�h����q�f��Y�sJ��P%���|�48W"���秣
����>��r��H'����?D�����~���Hӑ�;�F�i�|8����,;n;�t}8�Q~�1��x�d�rB��b��1���exE󬎘�r��dՂ�+޲g�����\�%ӂS|�ƣ�*�q�p55'�p7Z�U*`@���H.
3C� ��+K�u�f)�V"�~nDH%yZ}�g)��F���{ӊI㊛��BgƉ���F����X�ɥ����`�:����I�ݨ3;��_�>�� ��"'1�Q��	���s���Wq�S"�b�믍Z
��h�Vq���"&��?	�|�.&RO;�6b8r�<r������5�Qt8�=3��wd���S쿈���#}s@�)�B���a��I�����2�烁��'8+��4׉��'6��L����!�!���g�s%��D��W�T^��4������g�sH��չoWS�ԩ�C|��6O��W;�Ѫ~?v�>:��(W��i�v%nt����5��t�^�e���/���ǎ�H�!�a��lJN9��������o��%��Z�V�2��`#�8�����.
�/�0q
��`{V=W��X��Ț��>��C�q�4�z=/�fX{*27����u"TM@������J����t�%�����v�'P�Ru��p�~�e1�ٗ�x�8Ќ�����"'�N��5� x��e]i frj������w!�H�C�ȶ��iʮ������K͵�8k�\���(�LCV
��|M>=�}��d���"L��X9�2�RY&�&�ˈ�d��B@I�?�EzGA�ʳx�⻴��]�=F�`���7i&�u؋�����Sv���n�Ѣ�W���V���޵¦��C�0�UG�s��o�d(W-&��xs����{�o؏iͽ-Řc�a�6�	h�c�Uޑ�5[��5^���$φi�/�yvOb�i���;�F]1UX��֣H�>A¢n������%h��6�Ap◼�X��
��L;R�KL[�e�2�Ԗ�(�c.���F̩`���z�Z���.I0~�H=F�S���N`m��k�;�eZ[����ּr�b�J� �%�i��_�Y��=��'J���d����*E���3�]�Y]��mi�i�@(� ~,|t�\�N5�$��:8�}�V�̈́O}�8^s._���B)܄*�f`6vw�?����S瞰
�7�PIVkCk�{x�����O�u���n̴������?�1����IA�y5��b9���%;w�@}t�Q���w������Q�$�a��{ݞ������Ly��l(j�RrT�p�Q�U��`n�M
�Y��ڇU0M��2�ap���,0��4�8�B��Z~��L
���!���*i���b��ڒ�:�P����ELj?�  V���%d>�_���m�>s�)a�)�y�}�fH���r�k��)׋��5�ŵ�*�aY`�,�{1�T�a�J�R�D�y��~`�����Pr���`+h��g���J%�L'�6���H|^&g�"�p%���.��KF�Z;��1�������Y$}��.P�7XH<��"�u�����:����>�&d�Þ>�\����K=?���"�ݑ��6�k��I(�p���i):g�H���*����O�������˔��<���|X���9��ڮ�:�M3�<�	[&0rN��?L�A�Y{މ��OȾP�b�9&8��������)��`K������;���O�����煴^�_�~97 ��b.n�&���S����,c{����v��	T3m���*z¿��V�$Is@q�{�R*	1�����5�eJb�wG���K�P-6�?�D��f'��=�8�'�%͋
� �������ǍLv�瓈ȟ�����ȈE3U}�������M����AJ2δZX�o��+B�W������A!Yu����X��~����{�R�w�D�H<���CC�3�%ޫ�mU�{��Ʊ��q2v�eD�9�Cj���ЫZ���e���?�o���J�HI���4�h�~�÷p1]����i��rM��2] fB���#�tU�{�+uyd�y�l�hީo�6}:n%�aH��Nn�����n��f��FU��y�����0v=������鲚�8��঩����I����i�i����� �5��ׅs@&�v�/]�u�U�Ԓ��=���"m#�ӂ��X��ی����s� �Q�����Oh��'�I}��>$�~��U�臡��/�PS�5D��e8�I�z��/�86GK��1,�g���0��+��cu1�n7@7n�r�x�f��Tߖl�i��g��U�>
/�#��������YBJ��`�`{IaZaď.|~�k���ɏqh���O�;��_��ݺ�W��Y�wƛ%���N�x�=�O�
���j�ͥ��h�⇟�N�)/�K���;" $Dy��O�µM�>�� [�I�v�ןT��G�����;�*���oU��:(����:�a�s#�c�t���������ߔq��â�-?M���q�X��HrI�@����8��7�a5�um�u����ȾqXI�8Z��s����d���۸� j~����Z�IG�_(��̃�"����w��g,�NE��]�6n3�uD�����n]�K��=�9
:�:2p�<]
�3nƧ���B��L[�ՍZ�����m|4@��qv/�f�m���̾����UoJ��~�q�!���z����"w��L�����+��m$�݀xnd��r��c��%ݔ,p��3���8~i<��E �����9zu�B,���\%�}�9[�˕���9�'�\�Ѻ���_b�R����4W���w�,S*q��L�t?�K�P"����fƿ;���y�A2.��K�	�*)P	�f��dO���kz�3�J�����b�FGXN�5�f�}8T>.Ʊ����B}�q�z��ي N�:�7�&������h��z;�0**�bs �.��g�Z�I���=�H�wb�~T�����X��X����w�C��fofz�[R	৪{��ɠc�Ġޑ�0�2/��}�L�@��Q:�lcV�Y !��NO~�AW@�{1����#N/d�d���-����r%�<n�f���Ʋ����W̶�Pr�w�@�0I��G�����6q5q��ϯq�;%";Y|SlI���=D���;���j8��K����1 ��5|�X+�[�űv�cG�f2�6s��F��-������˫��&�U~� K.&-�]������q�{S���^��L�
�����2P##öi�=mVw��{oj���z�0P��N�r�����\�Е-������{V�@k�<��FG�ʰ����}�rUl��<�}�p<����L1<�V���������GpA���-Y�e�(��1n0�Z���u8�!�r�E��P#��4���������`;׹��n��Cd�������o�WE�dV����T���n]��T ��I����
Y�an%�sDܒ���
8
��&jGH`Ke�WHg��RL���Әe 0�5�3�VN/(9 ��4��~���Ƴ6�L�0"����)���	�����R��婪��L�����LK��fr�q�0�>���7YX�x�b�ڡa�g�%�_һ���o��\�8:�ͥ�+S�[gy��?]t�t������\H��c�Z�Jq&��Kv�g���<.�e�E~���۝�ңz)���u����Y��?S��f)ҍ���R�X���Qol�p��IyL�҅�%�Eޞ���WHs�b�s�J��h嘑�T�%�
{s�6�*I�Ў�恀�@��U�X�x�Q��)��l�e�׉,]�j������o�3�6L���W!��%����� ���xes� �R�&Ub�R�.���8}���6]n/���S$
dW���T�݃�^rB^Jm��+<H{>�c����yѫ�c	r/�U[�;n�+=���Q�K��a� *���#�!_�!�g��E&���*��ƨ�������fݕ������v�H.�+�Č�tKQW8�n�C#��f��!T/�� ��������-2)}��:�~	��t��iP���L���k:8��3�,�r{KD7
$�n|C��+ۃ=Rd��)�oo1�����Ӥ��U�{�n΂-wvKs(�rlo����0mD�#��6ٽ�T}��f!��4��0�F�$2�Տ��A��DP%UP�=1>(����1���?��/sc��qI�̹s��I�7�t8��"��e�TRo�lp�m�o�^U��RT.ͷ!�7u�4����
�ѡe��\^�TD��g#Doh˷�B4���r�i¨p�~�Sd��<�� �\@Nşpj&��qJ�@uC�Z��SVh+sw��a�t���B���d�ၭ)(�3(���
��% ����Aik����E �(�/6g���F A��	�Ĕ^g��k �£W_�)�e����&�:=���i	t²��+��/�R]f!>�"Ʋ�b�$��%ςn>���AuO���A;����j/k�&$��|�$�٤��X~Q/�r`֣�*_�8C�~��� ��̪t�Ƴ'��c|B0��,&���Ǌ7jH8��@���n�l�pb�R��M�j@��ۿ�ɮEPG�BQ��7�Be
~�nE1��M�#�9�� �(�� �{��|�������h�N�\��hi��+gs�P�^�6 ���W����*�h�br�����3�M&QC�U�+f9�p,[�{:�z�j��]�b������>ZKw�E�<=*�`'0�S�5������́b*x�m���]�9 �r����p������C���c>��1�1
`��!Ac1B'bb���r���'���-g��ǼQV��� ��x͟�
��$�uv�/`Ǐ{L=V��xp�N���1a@k���fm�=-T�v�"AC�W:��@��H�u�@\�:� ��s�(�uJ<[���0K#X���Q�I�2dw��5]��h�]t����`�]Ij]��Ԣ�	���D�.<�؅���F�+�'�n.i���?I�o�%��JD��p$�*CZ`�Z'vU r	C�/O4RZ�A�{\b"
��_	���� Yӫ��y���$�c�Ӝ�9�d���u�����*�Q"�����-q� �*�1u�}XC���e|й��Vv��UG����*���p��a�⺥n����Ǵ�a��
���,���M)��Dr/�� ��0Aԥ�f�YM��u]�G�k�#�D֒��(T)sOߴ�I}��/�b�y]~�Z@3�Wi��~���;N���f�m!��O0����DJ �z����D_v�񢧿 [^~����+���Ԡ�>Y���뷥�S���I�5����5p����d*���#�/�c:f(Wz$���I-�gH�j�y�d����Oڲ��[�FZ�YI�>G��R!M��]�P9S�	MnE*�=��_[ی����Y��/ec�?����n���#n_������`UR�xQ�OxjⰍ��6��+lUY �[ʛ ��7/����X�ܗw�>d"\��5�i�7 ��NN��hC����Oi�?K52�S�P�P�K
��_�������I���Xd͌��iO%ƾ_�������y��yӹ�v����Y��izN�.�zV��w�/Z�2$�̆M��-u&+5nLx�|1�Bط�4ud�,x�$1]<����9姓��^)wr'����[_�ߡ���ܩ��UP��͂A�UR	:��o��Z�ϩzd�'5Zzt^Eߎ��g�äH��R���8��#����^�L�v�?�.�̉	S�o�Ŗ��~����[8�f��#���ć��&����u��k�3]ʕ*O4�[y�E�T]`2��qm�)�6��}�
Ƹ�}|�^��[��K��C��D�Yx�:2qZ�
��*�I�B�
!l�64&���(���v���m_��Ef��5���NM�=)���	�d>D���6F'Hz�bw���wș��m�P����#���J���}��`=2�t�#Ȑ��;�N�U��ʹj:� ���o���
|п�;Pg3���h i�#j�"�*ٺ�m���*� ��;�b���%��'��c�=�z��j�8����
�=�nQ��fʕ���+!7�`��`����#b�cl�)�|�(��F:�1�O#n�6�%[1�
F�W�p��aޗ9O�g�f���0~�Tm�X���f2��o���C9��qmO��=\R����n[pt�?�0^�_��N��b�4mu���:�O�/�nbk�e[��Y�<VCҧi�À���/�	Ft��Q���&��\}�qr��}�U]6�(Y)[=;ga���I�VD��\��*�3̣e�qٱ�G���;*�ˬF]���8k ϙ�����t9k�"�������ش+A�8�m����%lD�z��o�|�gj�}6`�.Ѓ?	��C�����)� �"-�?�Dy��;�H��-J�dɳ��9�ea��`N^�)�dq`u�u�X��|^b�V�%
���������R�%ø6p0���{D�~$�T������������Tw2a0]�P�3B%��t!h7��K�,7���V��u���\�NXf���o�0���h=��V�hϛ�oڊ�Vu�WS�-����Cz�s|����qu���n�ߺD���P��@�ʏ����(#/d��{-��rI#y���w|�$�#o^h��2��叞$��V#Х��)�j�) �"pƜ���h��&\Um��F��aP/��I��,�@)i�T�p�E햮;N�tL�����?"�q��fq�g�Z��� �@d�d1K�Smg�9�P�,�HkŴK���`�Vn�X��l��M�U��Q֪��څXհ�G#�B_��V�@��xq��4�`��k�I����@��ߘu�I3�/�
��� ړ�e�xwq<X�/�%��X6ؔ�g��r⠗G�p�?M~�~���lvp����p��p�5�j����ߒa�m4Gh���ǯ���\����k����^�Bߜ�P��lg���P��r/<�~:J@,硾��s�c8O��ݷ���oK���_E�Wrߌ��Kk�6.
ab���@"|����,�$�\$����.�Q�l�WYA<��<�vo$N�ޝ�'�ըb��U���#�B�ox�q%��)^?=H�_ƴ�b�g��%Ղ�:�C���)� **�s5<Ѳ�ҺQ�n�1�j�n����-Q34�sG�D
���r>�nɜ�H�Ƣe�����2G�J�<�&�\��O�w�AE�)n�-//s1�5��)c��p�{uW�<��έ*0q�`��G$��qVO ���5�1b��d>R��ܦ��3�c����@�:`�\ �#��iD�MR��Rk���Y��������fx)�� 5���N�0xފW��:�L���F����od�C�$d*�H�����h���iv��"�ʚ�x��-�L҆:�ՠ��w�%���8$"-u�3
8�Y@�K`�9�Et�nDq	e.���$ �2���eV6g|��������ܷ�4��� oYw��@�]&eݪKS��z9�ڰ�N�C�'[f���q�;�s�U��*xk�PW�օnz�|�[w��g����xBwL:Ϥ�g�hV�:�)?��c̓j��a��%/��t3�,O��(�-���uw�Ͷ��X�%���P!$�v�'��q>���F��4�D���
["˂Y���k�1��eÜ�����4���ֱ4]��s��[���թ�Aį��]o�;x��^���iy;�!� �BS�V$�0���4Sj�̊}z��M����Ad�f>D�2���w�6�.Y{l֌��W������j�� �YyY�$���Nt��� v���_�x���7\�ڡ��c~�P�O�Bq�@Fgj%��Q�3��9�	��G�r³YqV�D)�c��2:`%���YH���]�����´���'�W3Y]��s���f��X'  �X	������M8���ő�8OMT"fw�k��)��0�*]UU��q���p�`v����O![��I�dN�h(p>��v���AS\��e6��f���Qb�#�JMj*x��E��5!ZaZ���̛���TR�c"�Qru�'U+���``�:�����d4�*�5��$r=(�?A��(�?�QP_�,ʎ�g: ����+1Dݞ�I��cŽJI�%c��QӢ"�&�\əxvo6ڇ:�������GwO���%T �Pd�|�؎�=�7�>������)�nsM\�(}$���� �e���݀�E_r5����c��%@?�4�0*g�J��b[��h��ŀy!�",��-��� �H�\�w�&k\��w��jx/s�t�?�
��̯��2z�:^%1c^=fO0|�#B)��
<Z˴m!27��Un�\?��G�-��|- 8�yq�z�G%m-�R!Z�ė�'���V'؜ �> �S�}�Y�㦖?�L
;���/4��CA��f�I`��)��oD�hȽWvh�Q�3�&t�G+jkV3i���~�rQ�,�U}2$n�p����w�]���Q��9_��� =6�\��olLEv6�;�C�u��B9q��'�?g�ñ�y�Z:ڹA?}lZ��5F��!���m�*)Y���T�ǵc#Pt	�ux;�T�����'`Jz���ԅi +�Am�	yk�Ĕ?����)���~jBѬ^k{��$�i�i�K�`�};��Z�B�p+#�0/+�B*?pr�a����Y���$��1����V�u�	��¡�Pյ}C�L�`��M|G�G�������_����<�qc/��g�-m�Q��Ĉ�R8^�����������c���/��Νi�+&�~q�S�ګ����2;��O��G�Z&���߮��(��.��에��t�&з����C랐[�F�d4�b]抣pf'��c.!��ȣ�3<<>u�R}�_�+A8�Kܕp��M���Ep%r���\��,�����8d�z]���<F6RѶ_#{즙��D� �
�SX���t�ӼS�
�?)�m?
�{��=Lo�������Y��@���^��k�|�����ذ}���X[xl�F����E�<�OM��ΥqI0��B.}iA�?`����;�����B|ޭo�e�1�-��c���5���Ѥ�e�Zp|!Bj��ݮ���K$�iVi�a��p5�Rʈ�v��%8.2��V�ۯM����xQ�^��O�2��&`�n
�jsp1��-xs�P���P�/tм�N�\{�=�yޖ`�Mq��\~V�E2f5�OZ��&5��%�^&t"�Ej��IV9�d+N���+ƃ�d		�J�ʊ
�6�{K�ˤ��X���Zl.��"T�3��J�#�l;^(ǫͲn9�7||����P���V�J�^��!<^�V���	0B���&�F\���zǕ��J�l}�Nv����ƌ�՛��®+�p���e0�V�D-���[Ti<p�h;C�c�q����*�GS얲{����+N]�s�]�fω���m��t��7��·)��G�ic!M��q#H^����#m��}:����9�9��7F���M��
��<E�z�������pψ�ij�K���<��g~%���*��^N-3@���vg��=����#�[LқD���$��s�r���Vh���x�\�}Ӷ4�����}�ʴ�|�;�<��w����Ե;�R��hC���O�t+�=��.!vCW��
�oD��X���~��h�dޘ�i<��|�[3y�wo�ߜ��7�^���s�螉�����&�T �w���R��T7�:)Xb�U/�/@D$��+��������ɯ��͓-)p�gu8�^6J��ui�����i�z�{{X�y�D��46�����ƺ	�9ې����3�&ǯ�"�p����/T.>v[���\r�te��>(ӗ�����H�Tއ���[��?�ޢ��x��_դ�����=���e2�Ӕc���aZ�e��§��ùK4cDy�Ijj� /�?!�������O�=�Ù۱*r�r�`m54#������&���%��D���u�yy�Ik��*Z&l���f����X���X抱�J7ᕎKU�D��ړ+�pi�a�����΢ �*
�M"sS�ZR�Oa޷�PC��b��]|9��Èfj��'?I�ʇx�(d�-�Z'�e�Q�H(x��B�M*�y��ͷ�µ-�v�ɚ�8�I۬$r������.�H����{� ��a�9��[�%L�*搰B��h.�lA1��y�K$U�B����L^�2�ϸV0�ٞ�_�@���Q���^����;9%3Y�Q��n��A4��^����N�7��IP-Jg�R�Nh�JGb�1�<��ZQ�#wY98g��x�4u�'Vp���H����'��\Cʘ(��I�:�P�0��ќ�5���YX��GN͎ł�':�m��i��D�,(8����Q�i�>�ۗ�7���q���2��Ss�&k�۴��9��e_��=��*���;��~�dg9�}[�H�G�G��)�M�v<[�®�W��y��V]����&<�f�
����,�g��I�x�#�S���{���7�����--�XF a���[�Z�e�Y�&����H�u)�%�
ך����-?���x}\�t�:�5�Y��^�R0���7�� ��1VW- xa<�ݓoĮ�}n��J=5S�i��r�YN��@��2��(#-U���YTTI��Cܬ��'�&ϰU+c�n�]�:��,*�aQ����e��^��eP'����u+�qS���υkH9'�D�5-2GdB�Rd�P�X��xٿ�!dl
%X���"���/\N|�����8J�h��L�}��_G�!ǻ)��\u�Vޱ�x�]��ݐ��,BD9:�J�3����F�p-��x���hj�-U�|�c�o;�L�ѓ��98��V$�.���bJ�c
˂�Dh�A�L��
��ߒ�n}��D����`W���#��G�A�i���m���d�a  �^ǀ*�I��ϧN��-�}h\�m �񸅍�@[�O�#�HLje>d�Y���Q|�^�P��}F�wt}R�Z�thw�|�$�x K�J�_��81]򛋊 ��~j�C�WT{�k��)���/g�����[�i(��8���?�p1)  +_��}��~N'i�xV�	WP���Ti)N��:��YD\	΅�aY��s�\��ϔ��;�٤t~�X�~:�f��rm+�|P������x���O�OG�HR�5�(~ʂ�L��4�ay���|<+��g�M0��NZ�X�m���Q�� ����0M���K>�� �d�B-�V�����mP����23�!�=mШ��j�_[��R��\��?T���/H�>]ty}`��o�淖�{_�:�c�˭��L� ;
�{"y��1���#�#���qT`�&V���ز��-��鱒�}�,�+u
�@I�R�ZNiK�csW~~I�~�s�ɥ�t���#sV�Қɺ!���ؔY�*+��o���+}9���볍�R�I�,�<��ט_�S"2�&:�-/ۇ��t��E�H�v��s[��21��Z�8�A�r�+8o��JABru���5I���PĞ���, #�+V5�F��KE�B+g� �G�,�)s��B�o��f��(|����=��(���ſV�HB$�SNzG��E��y1{��U�ɟZ��5�2DEa�8����nQn�X#�������\,͘8�zF{nFRD#��Z����e$�]X#rh�U�О�A'e�����'GPƶP��_%�m\�!+�!,���c�b�>IfMx��ׯd����u�a{�`Ld����kL�'F%p��1Mn`�Z�Ϊ����w�� ��sk�޼jwæ�U{wf��3�_���iZZ�~�vN�š֒6>�4���R�f^����T�3�0G�w�f�h�C�q�f��e+�Α�kE��w��֩� ��F~���9j�!���@EB�z�P��;E��L*7I%)2iN�.ׯXI�~1Q���28X�]s�E��J���A.�#�a��O1.:&��EQ"S-5Nh��@a�Rx��^���3�0i^�]�뀆c��f�)}3�b�f�h�H�c9g��P�k68ڈI�G�G�~��ʇ?"�
K��W�"j쯙\o@h*?����K
�'�Cy����	r���+����3k>�g��@U�yN>�ل�� ���v<�c����X�ZP��bkM�,��;<�?�Y��l'D	�].jA.W���ڒF�����IW�<�x�/��c�Ms�9��#�8GgG��Q$aޛ���E�����`-������wOO�S�����I+�d���v��ЙR.��H�)��%ne������Lo�G�8Xy�
��K�x�ǹ$��<��v�h�yw�O���?�T���~��+pÃ`���4~n�\PZ�+9;{tVC��I����A
��0����z�7v���ϥM�QxzI�)c[�S��Q����>�}ԝ4n�����z���bh#����UѳR&t�#*Ѯ���N�/�!7�n���X���N	oOw�,���d'BN���0�q���+�sU�|��`q.�8����)�B^)o��h���
�Z��ez��=�*�П<S��G�ho/��z�櫆�i��P�ϔ[�����7h���`M9䥘��r��O?wʋ
��f�>Z�q��L���p�si|��p� M�����/ĤKcN�����m^3yVI���������=�A i�@\�oB�]�X"zG�A��k����G���'W��8.�@�X�6gm�����%E��#"iSY|u5��.���s��&�׊����W[��+��b'sc��N\7�����]E�_�"f���P�����&�y���n,���%�0�{jm��IŜ�x;g`�Y�{%G�̧]~���#�}<�*�R|�B�a~}W[b�a3g�t@��2C��舝Jq�uvH���$f��\�O� �,��K�*&�.=�v����ht��:vs�
 U��͝�K,��v�ؕ���@8��1��9�z�x����+:�"Q��f�r�C�4�wau��h�[�0��'��`}�!`���MxC�����ǅ�Ծ��u�����dqڷ(��qE��Ht�"��H;��X���>.�g|��Z��=�������[e4���� �F�V
A)�V�D�UqS�_�Y�4F��J^�{B��=��A�;/�x�#�)���¯�8;��ܜ�{�u���M!�p��y�Q���%{��3�8)T�����դ;�ֺ�A}E�bR��)�S���DF'�7���]��V��I�P�%)E�[њ�E��~-�I#S@���P�/G_*'�O2,�5����Z��k�g�E��څ���=� S~�� ڟ�����8d�92�s�?��?�P��Tb"��Ŷ	#p^�Co6�����h/;B�}Ӳ�z!��6��='Y=2���>R�@q[��#�`)-��p� �oS
lPAg��&{��&����I����̞�w�@��{��a��}��,X�I�w7ƔPI��躋�6\��]���<|��p�G�9ō!���_S�/C�&&n�W-�f����咞�Z(x�� �'�$��w��eL���Ռm?�7��H	ui�iz\�8 ��;߱�@G'׼��\�n��=/�;c�T�#i�ڂ�R���vH{Y��M����ZsP���՞�C2�^�$�$��r��bH�::�O/�ڟ)"i���T��}U>?=tQV�`�H�|/�T�)m��C+��KAН���=�'�³iu�+�-<������J�g��{K��g~-p
�N�˪^�-��^H7�79b1��vU�ыA��&�rM��O�����NE���¨]U)�2[��@4�GC2�QH���h����i*��H8?'74�+^Rլܰ;o`��	�����/�WFǂ�aĠ�@� \�vk����d�!��>~B���

�UO�ёߥ%1g<�fiYB�[�'O�"9f=V&��ݕ��n^MX?M����z�9vc��U���ؙJ��?mAH2k��.E��&.��w��h��N���M��@�����I�]ĭ��i����/@��뽊��ZK����g!2T�,U,$���2W���"6��׍��-f�(�vʒ�w⤃���y��:���B�4��Szz|����$&��L�Q\��W����$�w���x ��R�B��:0JS���i�B#�L��]vǛ"R�@���,�*�^��|�$n���L*s�v������'@����СX<7��k���>�.w���3�̸�/@�7VHH�F�b�7#�9�a�������F$2��H˯�ٰx�y�c�F+^�Ҩ4���"C�̆��\���㏔��)Å�ަ@��_H�^����Q
7Գ?8Ur����<�\9�o��x����,j.ͼ�3��_���Ʒ7p6�N	���uKoc��1.�%��ݦ����n��qG�6�L��-��H,Ғt%	�-�&�i�w�H������gTCv&�����
�yXv�C�S=�y�Q��݃�3bR��a�=X���u�^��j|\���� ���W��Z��*C.��lA��Ͷ`�3����i�H����77�&U6�A�$��;��������FXΕ,f=5O��a����9Xjj�sk� 	�Xʗ�w¤�hg�����x�v�`�7�
,�@5Aj����΃���)�\f��fZ�o��t���Ā���V�m�>���/A�m�W��D����u��c�P������;��8-���q;�bd�E��\B�+��D����7h̓�lhb��-���+d�7��qY�>��
 �/ƥ�\�e�����s��[3 ��O���o[���{��f$g�G���w����]-����ىQ����%4���֥1B�A��|L͓��YʝQm��E�p���^G��YZoxlU�ӻ��m��n#$&�'6x3GCOn��R���������2���C�2j4SA��z�6���m�b����ټN4�U�Ҭ�
�8؅%�4���i)[>lE\a�lh�m3��|��gwi�$І�ٶ�,��ؑ1lV��R���XvvJ�9�URşK7��LF�q�I1�y�Wga�ZB�f��^��P�^aXvJ3>�S���!8UAqc@"@l�GoO3�f�h����y��yn�-׺���C�ѣ�t?)�=��g�tA��%��t떡�vt�4S^�L�k�I����E��_4��:��
c+74T[�c�_��W��\���SgN��IhRu/sX��hN���^��7��V?�eL�{Χo~q"�ވ�r�|�T
����8�DIAn�7S`�em���'��N�(mrP���v���dr�En�Sڒ(O�^
���mԀ�Z<��K�+m�$54��K�td��[0ī�?���g���H��>f����|�-ŢA&U$'ƹ��\�S�l�x�E��B �$��y 0ǥ`gw{�{�����[Z��bk�N�3�Kb��c�Gl�����{�N����?rC����"�,��[2^�Zy���"[*s��8:�nד^���/���x�r~�u�X���G���+şo"��#֛J��j���K{3��Yv���OT8�]�����IY����y$��7�*E��/6l�52��J� /�C�e��tT�܀ƾ$�Z����2t^]�
*���UO}TL�Gҹa��Ͱn�������W�]��h����S��k��N|¥)��_����o]~|�G�*h$	+ؾ��虾yS������W/����u6�lF���y9T{\�d��mk��Ҳ�0_���2�Ft4tb-R��R��!l*�����pO��e�q��法�tM�o�׹�tn`���G��=��f��#�I�]�9z��ub�:Cj;�ʎ��}����u+�(0w<?F�$<�	|��O�	��9s-���f.ۏ��'�y�zl:��Q��!{�t��7�hf?��C��gZ�X�=���~1�m����<���T��Ɵ��؞ ��wR@���k޷
�4Y��~��`o�x7}~��:��3����g#�e����5;��R���VZ-��e�J��p,�ػ��Y��2�F<�9�x=��<��i&t�o�=>sA��n�Nc`�M%��S~F�P^�t�)��Y���TQw��X,۔=�oa'����?g��X�H?GZ?\���Ô�uO_�hm��+P�g?�6�Mw�X���Ga��S�e%�K�]CRsvU��	�ޭ�\���(�d!�����M��(�6��v%�}7��oT2��=�^�q��Sj"����p\�FUPL!~����ԏ8�G�;�*z��n�F��SI�ə�s~�?���+��j��u��,h5ϵ����Ѭ�åQ$���d|=���oer�Wgm����>n�R�PDA���@��6+�Mw8A]�8�T�w|�	hC�S^k�'�|����L�װ���iw���BRڛ��z����a�.\4��`���
H�U�v�wGT�T�9�-m�O���4��
�EKR���--�p��E\%{�l������9�S�!�tt
��F(�`m�`>�gA�Hf�c�~5�6�Xh�ZM�l���cX�BʝS�3D��BY�r|��H��L��͑ޱ���?���'�Đ-&5�"�4�
��A�1�&�G�fZ�c�mM��$Y�Í@���>��ٮ�O�e�o�2��J�����ۀI��񤬟�hա�TD��F-�'��`Jb65��<�`p�T���A�#kK��k
.��2����3J��3J�w��ǰ{J��ҙ����1(������r�#t	7�3�����jdm�o~x��o�'/��H��Αϰ�2��K��k����WE��W#h=�������|P��`���:�̅G�XQg ؅h����ȡ���-�[��Qnڻ�~���
�hJ�l`D�<�v추���AL�������5,4/��M�\jX+���h�,�����	�:VO��s<�f���EX�܆k-r3Fd��1����f; N|�ZSNDv� ��su!�l��=����G<k�%�مm�j�w��3��p���S62Z�h��^C ���ݵ��*�#������z���Q���Z�ȃoHm�������OF�i]Z�6Q��
����8l(�6��m��ʔlݑ�^�6�6��!bQ�Y�O��+��βu�I�!D��G�љEj�Q��ڋ?��ھG LZG�K2�D^F��hB����_�#���Rj�,���|zN0xJM� ~�_��6�v8N�ve�Wp�j�T��͛J���Gsf\F
^z�|�&���Nw�qoG��x"T��!�VRu:������	ɠF,֔��+v�ö�l�n����:(A�d��Vuh=�/z��c03d�,��X�]D�lq�dJ�e7�)��0y� ۭ�2�9��O2&���4�<U��3���D���3�4m#B��?�)��%~���Ɛ����w�|�{��L��sʹNoKM���ë��Z�����gfϗ2��}��n?�`�_j��V����Q[��h	{ ��
���_�I����!P� ��k6u���1��t'�w�y�����'HZ_EO���wO�̅kѲ��r3<Q�7����d��x}�d-8D�HI��Y���2Ն�ت����6rT�\v)+H�'��7V�O�v�+g����z���i����o�8�S���*�a������ery�3MŽwl�[�b`�ō��G�%c��B�"Bf�3/4
�6��nj�S�3%=���6D��Hѿ�W-�b�R���d/ا�T�	���)�y�Li��h��I0AQAb܀���U�s>��V������ �?A0O^���`LsdU.��0lC
�$۹�O�u�#��i@�g� �tπ[��\���q��C3��`�Ⱥ��m_�| P(ѽ�W�ė��%�k�_�Uy��D���Ls��&��Y���	��`AY�}�z
���\���wj��AA�q]
�Qf�"c�-��5Ѝ�,��m�.S'�A`���)8Э(ɝ}awY\`�2�~������������U�/S?��g��̢��?[t�Wm_Ye�`�u4�TY˅aq~(�d��<[�"�.��}k������5wq��Q���KS�Z��ܫ�w&)Ԗ&_�f�K����w-ه�N�{9Y�%,z�q^�)�-�Kݬ���e�l�Q���qޭ�����WH�Uew9�6���UVQǯ*��c�|8�/�/W!ɷ���P��o����3v��J��,;��zH7ue:8@I��,.���x���6`�����_���zDY����ӏ�a�[EM���f�=�C�Bl_������i"ۥ-8��X�kU�~�gf��KxL�Xָ6�3�X�d�p	Fu��Z7�tk���S��=�3U�V���k}~��= R����Le²&o5�a�I؇3�g� ��WZ`s٘eK@ݲ����x�el�;�D�-��ځ!�쀤�R�`I��!�},�Yѹ��}����+՟�P&:y�z�T��&��^#��8jd���_�͵_>F�;\���K$��s1�5�f�~m�BH2�p��\��k@������w1�C��O�L�ڭH��-�PV���/Ȑ+����j�	�ڏn��4�1��G ?�:��E�B ���YZ�w�%gֿG�[n/J�ӓ���[�����T����t�����>zn�g��}�e-z�s{����`,�rü��^3�m)�/��s]��Wu��k�lه�F૓|c� �_[×r��/#$G tv#h�.�x�u�20���킊v~��������34���b2��4T��M���/b�Tr*qt��܎2q5,��溜Yhⴣ�
hd`Ҋ)H?aTc��b�����(�8��f�J��' �z��	b�n�G"w�"H��cxϛV�w��:�s?��
��H1�M��Vn�B��
�R�U|�����eVt�k�_Y��Пc�	�n�h�:�����H�ל�7;r�##�%��4� {!�<��m����SD�ƚ��N��)6�4[��(��\����6Y6𦒜�r��p�B~,�neE�YD l�x4��W��a��R7N���D�=z��o��\����<��z�g^�[� ;c�NW�zϿ�������a��}��9�,��w�/& �5���^��{qc��:�%��Z�[.�[vc�ºx���W��Qp[�w����L�T��y�G�|�0�dݢAj�w?�ʦ�[�΁\>��DH�n����U���0��>����2���F�	,�M��H"5�����0�N�y��On�B�Q6�袵I��?6�@9l�<��%[�+~(Į�m�1H��6����b�H��+B�D�T%~�O�Ւ��n�M��v����]�`1p�@sk5k	$�B�,�4�y����i���u��et�Ku��:�ݪ�ڋ�4��b26���W��Mhmm��X� ?�!��ʕ���
�G#��ł�s�WY���@���o�n����6Sة7��'���ȃ�~M�J�x���x�h����7�Q,B!�4h��*׻�ZX&	�^�0�R��&�����9y��jv&�ߣ�?S�
�X,�Ǥ��ek^��iD��C:�
���J���)���;yn'���LІbi�0�1�.�L�0�.�7��t;�a�g]�Ah[��k�J3�����FB� !�2ґ�ùx�'e&!U��+��E���ᩗ�.�A���-�L�����8�7��)���>�ޱb�h�'�~�v<�d�^�%��q}|����*�]}8Q�"vN���j ɔ�~�N��(%E'��3�*���v���S ?d���.�;W(� ����V�C4�Wcx�4� ��Ե�n����;xta*�:ieΩ�/`xtT�ui��?�n�z-`  &�dED�:{Nx6H�3��T��
f���m͐��,ܮ�o�h�a_�֪������MK�f'�Z=�ٹ��ce�|A�i/�-=�U��p���k���ʠV�uq4*���[��@#��.�8�`H�� z	j��Z�(�7��}�����x6�SM0-�=%���g�>���z�� ������e�&SEN�3�m��gS
���Y����h:��ؤ�&$�ԶYibHi$āE|l:F~֫��Y�����\)�6p�hN��S�\@mIz;$�b��<v��>�Z�N�*Ւ�@<b�5w������k�6�:��J8�M�ʎL@Y�-~?����2��zg�A)P�L�>I�o�p~/��l�>��+�:,">��'���c�I+���]���k��T����aZ�н��v�Y�,�6@VD�[on]�]ȟ������m-\cC�H���:H�P�ں ���q��;WIz	���wt�>9~���@�l��Uo�v�����?I�Ѧ~܂ y�}h;��	��ByM'�G2���'Ul��P�6��K���?�e{�;}�$G���ɒW*����Ƣ��2�}Qw��ځ~=�<Gr9^i߮�ǔ�u���o��|t�zA���od��3%~`�U{TL) _����T������o��R��H#��c������t�8��`�{|�� *ـ�B� u�?n::<+|�~Si^�n�zS_������O��k-�q$�D��G�v���i����qB΋�r;�"����tS��	1�p���`���;�6�ȞvM���!��-�������O�E��/��C�_�#�t�d�]����rd~����q$�o;5�>�gy[�
���e�ʜͅ�!�����6��o��B}�|IB?q;F���t�T�3��j���ߦՑ8?��_�v�YǙ��W����*���m����w>���C�\x�7�֑q�gk��EP�gz�Z�UQ��j�!]uR��d�CS�)����m��1��H�#���C�0d���9�H��݊fy�1�c8���(�?Rb6�*=�g���Rѽ���*�zu�@e-udx�����|��0X�f��(��X.>��gJ!I���Q�kru҃6�/�w�ZT�}��i�O�y(���V��e��o�(Ӎ���TS�Y�������������-)\�x.��KB���WI�2CY��rWT�e��K��l6��I�v��
�6����[����k���w�ψ�5�C����[��X��߸G@E3��rd)��ճs X�_� bۯ'��Kw��Ė�ͱ��AB��W�`��F׸d�a=YȭE�7�]���w���`�{=D!u����L@�W򧤁�gd�����4ى�x`[)�zi�D��h�Cɀx$YB��"(����;*��Z��~�Z�淚�*�{q9�&�s7�scX��<�̹� Ǖަi}>�U(fո!(g�Y\X�/�1 x9����i6��9)(��0�����J�2�={i<�,���cI��9���}lW{��;��~`��Ka��`��rgtR�`�%U�H��E(�,{�C��G�I��[�WO!���L�cǹō���sTB+PRb{��zxl�\�AкnDA[:����+�aÐ4��t��
����~�{I�h��V��ڸ$A�@dݳpt� ���M�%؂M��7В��9n�6%WlZH)J���G-/1�h��q�Z�C4N�Feg��C>��׃�=Fd2F8hs �����@H��Onɔ�ؽ���)Φ�Z�I�ap�d5���Ӓ!�k�$%z<��Oߤ4r�vdb��+xח�U	��X�&�d�cbm����&�I�%�յϚ�t2�	�����!�U��KQ�f�x�@ڸ����������S��2�yÝ;ޝ̍�2�҆	�[��l��jN�VQ�\u��OM�f��`=&�~�"^�<��`��ػ�
�i�/��:$�� @M�W�"0Ru���\-��_�Gl�rq�����KgN��3�F6%4�MBJ�{����9[�������
cR
����Hk��ْP'�1���I���+�T`Py��5,Wi�ض��i��7�ό䞔�Q_Mrሧ���z/�bݢ��g�[ˈ�t�?ǆ�����H/l^�x˳3�S�Y���1�Ō4�g�0/7�7�o�H-C2��!����WGԫv	1��,�L»�S:�����q�܍x�;��>n"uO��p�QL�gL+����S��W��z�f*>U,��͋���JF��E���I(�#f�AE/1�WSeL�Q���)��W��~�����h-�CP�/��Wus)RV�������N�Jk:"�`�h���s�RiZ��(G���$��aX{��΅pBNX���D��g\��ϥ�����E� Q�nh{[��4k�QD`'@>Zb��ܭ��HKB)A���1	�?Ӭ��w���Q&w��A�C��7�@6rp�F�^ Z� �O���v��Z���?��u �3��d�}�O�O�#!
W�]�����Ƿ�h��ӐY�	�����K���؃�h���|��]q9cj�u��N�V,\o���]9W�噣�*|����^~����4�c0���Z�B-V$�j�qQP�b�X�=>��_�:UJF��@8�LБ	��!I���3�Gd��>	���|ά��ƬÎ���q�~r�2X���JT�x�B�)��P=�Q!x�c�Up��<��O�mG ��(�
�I+���L��.l6ZO��6ѻ+�
��Vغ�]S�/=I�;C7�uro�R����S��ˡH�'5�G�:�(|hW0��_^=*zk�������s��:̛j�&��2�^#Z��A��DPKg�R��>��|�kQ4(ˤq3�Ծ�9G�Z%M�6�E\���֬�7�n ���l�ND��.���?ȼ��ٷ
�N\͞����rK��uƿ��/W_1��Z�����sc<�c����H�P��6<n����I6�@!�r2��]N}�i-;�T~j��"��C�c��ʙ�?E��v���C��� �`�<1O˒G��
*�"3^4��� ��1R�졁�#�n\ p�� �zWE��;�|��#R�[ǡ��(Q������P��ҍnŏ5g��W�U�*����[y�p��B�C�%���ljA���Y�/o���P�����Y����p7�Di��,#g*Y�����Up63�3��� ����Ќ�Ks;��R�I�} �8�oKI-���!%�l�m_��vJ���tW�m ���F�D��%u��#xx�xc�R�g{ERAI��#��X�����d������h�{���:������uJfn��HP��Ip�wZ���AT9T��𢋫���t��2����%K!��#��`�BwS8��U��bh�QႴ����;D��� �=x0��H������\��D�e�������=�T�����Q��αy����N����}+Ծ'�ӉD\	u	��ʯ����o��*��U2/���{N\p���J��E���:9�C�z�-f�"��l��B��|���w�(�anյ�1Yjy���͘��lR�i�����
_pE7Dͮ ��[�<d�����.�8r��ʄp�$����F�c"�n^�����K*97�E������
<7�s�?�vxq�/���iԧ�)�m_K4��˴�6��׌��M��sFU���˩��cB�4�2
�d��p��S�0t��8���܃i�Ob�-1,����N�TL=���mii��`��ON��9�ĦӐg{���`�%�+M5��J��䥾O�����.�XCɱ��S�ʋ�[�4��;ݵfc���E�J�2��3��6l���vl�Cf�#.�f[�0�^M�[�la���U�3��ҿ2��ٻ�ϴd��+�I���'�������^��K�@�[�]dd�s�r�zd;C�/�,U���E*�ǦVk׿���(��j�sI�h���;)�GaAo^��hi@�����IN_4��,���Q�)��1��eFۂ6����|�:��
�D�se;����守��@��C�z?핬�/�_���&�� |s��< ��u�k�Q����?��$h�l��x�A E�5%���g�ۮ{��S�or���r���"�RMJ:�(�;_{9ុF��,�� �͂o6��g��g?st�6�NF ӂ��g��3k���}�ɯ�f];X+�W6!���
���>�ZPRh�#��	�%���\�?ni���7�~L�^ �]�ce�Qy�B��;Gmn�7r24&!�;��*���ɼ�4�)�h�j�w��ތ�r�.�}PZ�EBE
��"�� ���/�K���~ϣ��9,��N
V�_�����K"�~���������JK�����b�b�eN�
L�/�e���Wͥ�\��h����u�1�u�d0R�m���ЧAU�j+�U~�o%���+�\�6�/t<���{����)�t��<"�� 
�݂��~ 	8_ ����� �]ц֢\�T}�}���=<��>�����"��/ܕ���E��*9���1��5wv�D�s�
d��w�����gE��ex�v��p�͋��tcI#.S�ۇ��3ؽ���p�on�sͿ���h��#ͤ���aL��mO�Jԋ�َ���2ԁq���L�{Ί����6R���J83!���g�l��"B!st�*�N��"xN?8-f�� �]���,C��j�ilS/F��X]V��q<&lȵ�]	��ӂJ��y�� ��?�e�/J\�!ph����!C���&�.����92�x��30���K_ҏ�QR�$���9�;J�5��vS�ox�EHBkQ�$���߮�26-�d,AU�v���З��k���>�u�20���5=y�q�3+i����\�<�n�/'M��n�s�|Nmx�Ǥq�R���k
+���d��b����z�zxq�T���j�Im��|j�E3�G\������|���g�DP��>��(�5�5���Rf��p�v��)K����ޯ�=&E\�����,z<�s`����$[1�֤���Ͼ�y�5�љ0A��&�W���5mXV��,��֭֨��~7�����Z� �4�;�����9�OPn�4M@����֗���7��N� �^�K�$.$7�*&�.�Ӏ��9	�nt�K�Q�<����s1������:%dc��EH:B_(�?�&�:������}�ٷ�Aa�b����5�.M�{'s]�x�9��l�F8 t$I���fO�v�R�k���S��}���R��^��- �8J��S&����"}eG���j{��%�J�")�J��
c #��[�3�(��n�`Z��I���k��=��i���?٠'d� q��Tú���of����$сo�خ����(�մPȉ��M)O�|v�RW���m�6�D�5�1إ�c��laOi֝��j���0��p��3]��I,U��aȸkk�~Q5u�ʴ�\�W[	�������ِg��'�Y�FQa%-p�]�GY��Ǯz� !�`5�����"3<��
ǣ�T��E?݂���a��G"�i�z�c�5�K>m�*� �d^jG�= NwP-Eۛ�Ipz��X�o�lgG��`܊�k����O���u����P���mT��N��,p����}%?��(�N&<9��p�K8��ͨ�\���5�І��Wˁ(�3N*��[�v/TW�^Y�����Ο���PA����7�i3j����1+�}`�{)&1W���I��i�������ͫ
�L��t(�4���{��w�p%A���1X��L���}犒�P�&��bd��fev�n6y`i�~�1v�Q�n�Y��䩇��3M�<��C8�	���V�w��ֻ�7�+f��v+�c�elkb6b{��7��CZ���6������W�.�#��6�s%t��Pq�D��t0x�/��T�}0��E��q����ȫ��_eU�S�l-7/�$���E�exζ���?��f:>t�*� ��}��=*�Mr���	=��>�%xsZ�K� �+�/,zg�c�y�z�d"sy!�����?߇��,Y+���	�P���؝�B��0u0X*7/j�3��Bɣ�<Ã��ŀLD�L|<c���P�$�+W��\4�:�ղ�8�OЯ̝��<�#�x����8����R9�5A5ˏ�3�(QQ(ܮ@6lӆd�� i���4œ���q�W�}qt@�gsj��b���ǣ�u1��
W��- ���vMn�yJ:.�����Y�~�c����f�8ZT�*��y��b/_q��yV-�u��GÒh���Ӑ/��x�wGȮ<�܁8�e�\:����}�3����!�h L�w��pS����dҨ����gK`�P�O�����q�'��(���8�2���5�>�3|$]�qDi��oX�n��q{aȼJ�K׳��vQ�I����Ӣ��붭��PbT�9ƒ�qY��IWVm�r���s���1��kb{,�������KD�),o�C���5� !�<�V�x饻��՘{��/M�տ��(	�>z��0Nxf�
x�P�#m�W���NH��·�8�$0�����s��܄�OSS��Q��̾�a�70�d�ĤE ϰ��B`�UI���P���I�R���p%pc}S�lrXX����h��X�B?5�i"fΏ%�=<A�jv#��D��%���f�]�ax۝[pMa�����ڱ"�[qí�G������/�B�,�fL�x�Z!&ai]��p7.+�H�n���4�w���r����P��JYߨ_�g[��xV�1�����yn��N<���ܽi�������u��F �2�^ʎ׊�}7=w֍�:q����ܨY���eu��c(]��S�Qt�J�F�
JQ�I����nh�^9�"Mо6��ϒ�'�c�V��\i���!	��+�Q~�y���,K�:������F�LI<V7V���x�����1�C_��L� ���g#�ǃ>&���J�'L��ߦ�����U���furi�4f��R]Olj���%3�(mK`I滪�A$ @f����K�f�0�Gt�p�۱����b������4h;t�̏��pz�B�������9�@'$��ﵵlXGt���ҡ{�$�E�7PW?�?��2*jI7>�� �3�i<1�;�Uv�.��7����]}��Q(ݪ�@⮳�Z���ۨ����@Ʀ��A8�9 e��^�'l��?P@���_Yp� �7�;�X��C�?nWF�<Z)V�6���Gv�����k���:�!�Ս©6pߝ�-��:WR\�>�Wp����P��+����H���:�&�k��8���kn�6������Z	�{kC�Vَ�����el�	c��C�+�ͥ�ߧ~�1�z�Y�F�ᡭ�5ƙ��{F�z_�N�"����I؟��i�W�??5o�Z�0������%G%�R>:�b�$C$W�E�Y"Д2�HFe|n��@�2��q�,��T"��lME�ި��gD73��|�]��:y,�/Z���	��yf�����|ۮf�[ڂ�9N���A l�町�;R�='���?@�H�QҶ��huL"�o_�9$_}&?��ض@ձ�,���Um�є?�2��O��m3K��^���(d�2Ǡ�p�x>�>Q+�J�7=Q�w�o�)���ě�߰�
	m�.�Y�ҳ���I`O�.blhۭ��1O�w�M�2�Y$�,�)��jH�l����J��� �q԰Q���̅��gJs��sґ�ؕ��߈�XQ���1���fD���w��j`��˯��ۦ6�z�RV^�oٓG�aj|ע�9ŌL�y�Y��FZQ)��XWck����x���Z��r���X^��z'�X��Ί �"hyH��/�%D�&l�kv�,��1���q@j:�f���]���(�V�ywoD6�X)��/�� �׶ႁ��g�E��
�For�n\��sVraY����ҡ�� b�`a�)�8n�-�5��~+�z�_o=u�����1&4ZA���P��z�p���"2J
���e
m��̒���o��6��ty�����D����(3ʜ��q�Z���?��ϩ�O�A6OD`�M@�jWu-J��ס!P����qe��H�����B@�zE"���k��ݏ���b<h10�%��s��E
�F���b
-
3���@��>�x���"ǜ�i�'8d�&%�y���눎�B�x�|s'��3���Β,�-T���%A��,������!i϶��>8i��<y4��0_����]}��S-�fi�fu<ʝGJ��\�},�Ӥ�K��ަ��ph�Տ���7K������n�$�jݸ��sJR�))��Dr���L**����	�8[?ǟ��Ʊ)����-9�=��s���
>�
wG��m=�,%�2�$I���}
�Ε�3��.-��T���UcN�$<]I i���I+}�sQ�G���"r�ۇ��zQiP�O��L�%Z�%��'�U>S�a�j1�� eG0��ҩ���-�:�"���� ��|V���	4��T o����d4�3�XR�,�u}�U���|��c�GB6��$����X��1�����?$:��^�f9T��Az��7�\af<oüս�t�&�U��CcU�B��D�(Ib�F��R�w�C�p��/�t��P)� ��$�(([�f��ƴ�.�ؗJ��b�Zf�Tim��|�2i�_����m�-$��dH�=�yB�cΨ�qow��0�9@������7�l���x�#2���V�۾��R_y4[��+���N?����9�CRy���w!�׏!u<o�B�1J:X#�@�Io0�Y�C�j�k�D�ldL��.2n�I��B�$\��)�U����U�x͉�rF�}��v��7�Rjr�yS^��*d�����%PK
����~�3p#�"�[���H����?�@'��o�����6fw��O�4�<b�	,�ЁYL�6���r����Q��S��[:Ў�9B�-xgS�D\P�13S�N%\@e�:���B�m�h���@�b}��nq+*6B�����V���v-�5�}
k�5�	%H�$��P���vrp���;�f����E���1�-�	؆�b���>C�D�q�T�ǯ��6*�#�&�n=]�,�v�/�G�9]
��t9��d��9����&�V*���d߂��.���r�M�S�"�yfVCc�	e|��d�9�����v���,��c� V���.�ca�#旰 ��Vm£k��-�K��{-=f2�:5��JN��n���Z����y���t��8}�1�*gS�c>�HD���/�F5�l|��$�z6�⦃��h.o����F��x%�;Q�+cAp��T~�ۖ_=�W�� �My�*ϝ�tJ��$ֆM��h^�ϐ�ĺ`�R�Dl0dk��qV���e"�>Үϑ["�WA(���w�Cj<h���ީɢ�N W�L��t���^�݀�'B<�����~���*6���K#�����R��Tx���\�lpzn�-�SK��m�4Hl'mG4!'�G�"8���w���ن��q�%� p���K��9lg�ql=�?r�c����A@��J���m� '���ꉥ��~�V��v�֎N������6_�CG��,Ήc�N�R�Ǎ{�4Ȯ^��������t�Wt�Q������nGG��ln?h��8⮱�Ђ�j���}_��"���FM_|E-K�%+(��F�f切=4yD&�2�p��[Ga��,��A�?��?T���&[�_e�aC�����q���5r�� 9�T��{���WT,L���1���˩w �[�5�[~�"B�5�pG�C��j�ԏ�$�L��鸓;
�̜0����Wm����j\,A��3�n��������ꥇΌ}�EY�%$T_�����׏���x}���P[8�{ 2���Tr�ڥvR�2�N�,�Q��1�5	ײ���>[;�sYu�ۉ��� �#�U�S��n�n�Z��k��X�p�牂�b�����:��h�.�� f�%�Pz�O�'6J�n���h�d��q'��m���j�8�4qF�{>�\��!ӊU@S_�)�ܸv�8��Rp�e�O6!
q
�v� w�F��7��T��R1�S~�X�(�,t�D��X�ݢ~3��Ȥ����o��)XO�ud�T�\�]�g���F��A-�/��Rs��i��W�
YI�wY��I��
Ŧ*?C�����\�e��+��u묟y奿��Ś�Y6��~�?��v��n�&:�dc��	q�韯�֡��}���	�άn��w�˚��|�I�C����r�Fw*9�?e��Cġ�u�Xc�t�g3�3���"���K�={ϑ������ Ә�ۍ���<��}En �3ы+_|��_��E�kdµQR�NS`��t[�6��	�H|4d�������ME @k�)�D�M��O��¿Z?��;5�s���8.Ry ��v����*�����or@�rܤ�o;ku8~��F��oP��[B���/�d0�����{W�!�DVJ����4��PD�{�ax k�񊏓�iO�I"�����������z��]�V��c���C.=yZ�Ч�ʂ*����G����j*<]2��3��uR���F�G�.���뜾��Q2G�\�ɒ)
:�Q������N��R�-�l��� W�����F�l=��P1���e�l>��*6�dcĠ��L��;���;ә>OL8W] ӡ��Z(jM�A�ST(_�VD�&!{ARx� ɻ#|����2���+�N��
!S�� ���Y$�.��HW��c#�{���ZT��'��l��;�*`iV����g���ދw����N�`�ū>�\Jc|r�1���FO��-��{�q��P����loN�Y�|4�C[��Lثco����N�K#������Qes��&S>5a.B<�RȒ��i�F�H ��>��\����	x�畊���u�Sc�CY��%�ޘG'�;;��l���6�7�9�&����0���rj����(�/���99|����M1x����Kc���D��9/^}r����ҳ�����j��y�h�K�`�\J��DO~r?J�����V9���Pʫ�����@Um`f���\`^ ��ڼi��w��4T�\	8g���?�$�Lļ(~���y�$J�;ф,�v�EkT�+�;��O/��cO˃�s�U� �ֿ��{l�c^+���m'���������a�����oeޛ6� �����uأR�=U�OV̿�7�p��W/pX��u�L:�Or�WD��βv����`^ �c�8�d�<&1�m���_��ұ}���|��HǽE�P��{�p�Y���ss�n#��%z9����3��ٮ���!Dc�H�z�j�y���[D{�R.Ҕ�庵񸉸��JT��M�I��σ�ᬛK"��0gHCW�CZEGApfK���=�AX~�Yn�&��dU.�,�#�w�����0�A$�{�w4+�]�.kyG��$L1K�bH,���U�E�yE!�h��Dp�Y��4�,�i��7:'��&��?1��<)�D{Y� a@p�6m�ȶ|�š����S��*ղ��Hni?�*�YZ�t���x 2�l* ������0�nr�hƋ�MD%���X�M�΄������	`y�?:)�0�O���"��7��,]�v����g.+ֹ�d߾�Y$&�F8%l ��p�nH��w�9��K�L�f9|�Q�ӊ��u'�UpJ����`�)��X6�Od��_��R�������ݩ��o�E)�
���&�R������X���%>�1���~B3m8y�g�+��۲�z
��b��,0���5�M|�,H�=��sQnP+���m��kH%�c��`��=[���قL��ȗ��$�A��_P����T��"j9��r��'1�Z$x�|����-�ցY��������������g��[XxFq�$�U����҆�`��^:��cq�����j�+m�Rcs����M�x"\ X:�^VGgh��z��	\��4��6�G��rA�G���"���tE����~%�H ��; �'��𸀪�獈��u���/���j_��}))k�?lz�;�1U���� ������CT��i�f]�.s}?�L���\EwU2��'?X��Hc�ď7�Ͽ%����~�"m������5�Rp���)K���s>�m�3`r����6�憣濎d�����AW� P��c|�&�ݖ����a�! �ʸSY}�x�v���R�j��������@&��B�����(7�ܝ`�J ���D��5zXhc�H5���I�70���YI.�8ʝ���ԋ��t>s.*h�c�Eߌ�lv5�L��IO�4Pj�T�*y��|n[�b7��2Tn��j��?�$��	^��<5��LK���[j&+���M���(.��I�oI�=�U�O�Y�UrG�:�j�Bs��B&�M��%֭�]@��_%������"1��-O�S-�`�Of�=S�ûn?��	�/����;����>�i��\_��%����B;ңfۖ���� B5��Vj�5����ZAj��
&�"ă����s�������~��Or�3��8@����&�Ý֭��w-K�?=�P�x����i;�xe�Bn�;O�e>��R$��}Ft�����X��._�S9�����ef-eJ�0��		o��P16!�v3�d�e��> 1�����BY,����.��PYtY��ԽY�Xj�=|�d��,�����1��&�s�66��֬�����n�;�4 �7�O���ú��J�=�܇���\��8�����s�!��||}�8��H�ɋ�A�tVS�d��G�C �V�~�~R�[	S�z`7��7��ʎ��ޒ|%�n�������H�I��ҹ�_�b8�뇔���rЕy�k��s+o�EZ.W�y����ؚ�j��0��HϨ� �J��v3j4�L"-��t鿽aT@� b���sڨ�Lg���*[>d�/p�;[8t���3�o�� �����=93�Zs �����~��`� ��zQMӹ��-Y5��7LQEX0sB͗��>f�h~UL�G��>�z�"���&�����S�.��.��0�%Owo�Y��Z[�Ƞ��/C�FK��ӹ��b;��x�7?S�/G��{������s���|�n4��ǘF��Gm�*�S��� E��2n�iS|��7�j��[S�p�I���2"�<��6w��-AX:/��' JͮsN��kH��5G�k|
��>s��o8[��Щ����7h���6�:I�/��E�P��rL�X�<�4�'����G{_x�uq�����`����z�S���m��Y�?/t���*'�������+�m�6���w^�tY�GE����.�՘N�k�;��ٵa} ����xټ�#̩\��l4{¶\ɱ�K�V�����*DP��ݣ�k����vt'B��˺�w�I�G Yv�Q��	�zǡ��31`��&�S�3/�qĒ���:���m�[�lP�-X�E����k{
֢�⏧CK�)���n+��[lV��P��T9��|>�n�������ͮ���j�V��5!k�;��G�~,E1�j���؆���FUxևj	�bŵ�x��p#�?�p:����)F_ŗ�L�#���>�dWm��z��0��:D&e皱�U��V��4��0�U�J���n8�(���+���"��fMnQt& ����=}���M����:�G�l-�{PV&B7��]�?�6{f������n20F`�֋?M�^�x����;�"�I����$х���f^^Yw�s�>�~�ڳ�2$UF��BVlo��9��`�>Z_����+:%½�~J����?���F���O�<�^Pև;�5W�\�1���:��Q��,���WqbM,��E�M�I��i�:�l66��1U^��J�V��'�ŜO�c����m��I��)���ߨ��p��� ��x�ؔ����H�{�"�
�o����n��O&��e��^���;9-�%k�:'��0���}�8���F.�/��U�1:z ��O}®N��S��אͺ��-���
6����#H�\�9r|��� jlu���d��:h�Q��aKL���`%�
7�d��3�������0z}����_�eK���h#`r%ju �Ň|�"��
��K���'!��V���W���<*c:�t���>�l�_�v���7F�$�mO7b���0m�]���뒲����T�r[c_rG���^If����_�nU��u�Q,�mo�J^��������^߄�ۂsb�_z���������h�'���b����J���\V��v}E���K{��}ۥ?�}��/�\ƨ
G��Sz�a��[�ۚ��S�X�^ݱ��D �	{��>E�x���G�H�aän��c���П��y�� Vv��i�r\v��+�/�}1/�2��*�6�o��d"���6 �ø|r����Z.�TO$�9z�M�r@��$��L"+\�%nq��2��`g�={�b,��خ3E�!����Q:�
�e������2k
4 �@������nh���cs���J<�b1�p�\�!�uF5��l���Nlļbu�3o����GÄ�GlL���DK��	��ď�!���?�����Z26&�#7|�����Z����s0V�US2�b�?�Z�l֤��۽�����2����1���1���	��'{����Q��\CLΛZ*=^5U�ӟ�Ļ�ޞ�CU���VB�u�,U��@��ki+�?�iM7+L�{}ktߜuBjӈ�z�GD�����q�zT�B\��-P^#��DO��И.���x-�#�ڧ�Êvfv��7��U������Sv�\28C���;�"����/_4�+>�;S�G�$��;�Z�s��ҽ1� D�_�����YEd4Zua�+����'�1�y�U�i�x/�؄��v�p$9���~���I��Yc��J��96C�""�͙��ΤK:���b��,F���6�<�k�Rt��tuE�eHF�T�>э�����`;(���3�g�ee9d8��- )���9��z(Y,��- '�~���S���V+�b�����褠@���V��6����8!��\V*:�:��r�K���'\(��Y�եq�+�l���G,����-�ߠ	y��>i΀�FSS��0D����)~A�s��r-��9�0qhO��PB��Tz�wз�?$K����岾[�KxZ�����{�����/���]I��5��s/�E�䮂�/�8I,EV�D\�)P�9�K�Ψi�|\_��:�?id �&n�]!`�ZZA���+Ӟi�5xH����|��2���ȓ�`�zͤ/c���bY�w��G�գ.o�r��j_�X���h�p����u�9�"��T���VH���X���@��v��IV<�N�]�����Dt��#Äx>�_�:8dS�-��]5=���#|���NA�b�djà��A�ܥ�Rj�>��Ӏ d�jH��� �6�Ƭ���vƳ}��E�4��G%\Ğ�*@�ݚ��+uK+l���j�D��,I8t��ZwcS�l��,���U"�11�����n?�@�|𚨪D�h�R3u(H�[k��bZC\�	F�t�:�K/6\��r@�27��\�� �ֳ],x����*���2�$>��x/�[v��@�9����f��d�89�%�hd�ً��!�B�e֥x�~о�P����x[;|=q5J`!�;�ؠz;;���4_�o�T��K�Z�-�rE��c���&�uhÿ.s-�u�ǁ4pU��׵ZS�����mY���k(^�A��� ���ױ���*�$S/�z-�d�U��A�.�7H۵�w+D�e/yʉ�;�/��Pe������&�e�����J�4U�{;}��cMϝtŞ3�x��<�tkF雏Sv����价^n�=T�C���o���5v���á��Z�$�|ч~�(։Eg���r��A�N���o�p�=�	O����`z���K���uB���`6����el���ҕ�����:1���!]����vK��C=�#%�Smw���.7R�kR5^�G���a�mt&���*;߸����=*��@̓�-g��u1��tqc�9�@.�.e��3M��Fr~*����n��_}2*�^Γ��|�|N�J��8����JMA�mv!3�Z� ޔ�����^l�N���6]��{Pl
rc܊t������!A�c,�x�\�D�K �r_�G5⹄�a���OJ�-��#&�����y?g ڒ�q٬��b����T	����2w�7�>P"$��m��������l��l	*��!��S��֞�_N���.���d���T��ݝ�P~�*���G.����9��0b0+�L�z�W8)>��T˨�Yt�>>�q5YϷ�br�/0g�-/�~���WkJ=(G:fB�~��X;n,�"d�$�P窞i�"=��T ?�Io��h�����&�.�	���=A�RǉH�D�"$$�W	x!^j�\kFB�5 &ܼ?�,!�4�E��*���R�L�#�d36S�3u�&�[��Q���A/[���u�3gZM��p�n'�������[_}�G!�!03E_5ֿ��=�i�L�u�h⢿��������R�b� x�3�&(�"�g��5[�������Sa�5��E�r�ht�5y��-�׏U��#�gs$�Ձ�N�}����ix͏�E�r��m,����M����\6ir�����\��=h̗���5�b]��mA��I77���;�e���V�5��8F<\�+ym�V\o��h�}+4��B�e�X���`&T���9'��0�0Y�$�'�
�����n�����'+@�lݤys�r�K�c���Q���P��1���ܼ�`ß��kS��l�"z�h# Ft&
� ���rnsU
��[��_�Kc�n����%i�	u<~���<�;�6����Ջ�R��'判F��MF�%��f�$vɳ`S_���/g1RE���y���l�]v"U_ʙ�hVbb��Z�2��Ȗ{�q�P0F/Yw��Y�.NJ�.����o��8�1fA���DR�7o���+� I��a��{)tr^萛x�*�zΛ��+`/ρu�}�D�=�OD�9y�ae�w�YX&Q�8Y���jd��e�ym����`�s�����|���a� ˤUYx��z��~�zl>��';���Gjr���_I�s�"PF���2�rF�*�d�	�n�U�����{*�N�]+�2袹�U��	�`�5nLR!\M����y������TB������)�Wh���_��d"Y|S��$[27���F	x��8�=*�S��>KXJk LԔNJ=}+|����%���Ɏ>��d�U.²(j6p&z�'n��G%��� �ٶ	��J�{gs6�y��ޓ�pZ���2$�����(>=_���4�z����
�:�-���}���2R+x{;��
���6	�[�JwJD�]ר�|�Q�d�Z�k���m%a�.�易��I�I ��5�5݆��]��A��y4tU쁆�x��u$b�n�	i��
�28wG��o��l�3���pag�v"�"�3P����@��l:n�'L�������3Lsn�Bt�e���x-�Z,~+�GI| �6k6><�g�� ��X�b�������6�h3�P�*瞽�Kcޒ�Â�;�,A�א9]��M}�J9�H� sR�K��֭S\�#X�����]����9�d&��2*EO�� �Tf���z�E�Sin��+�Sz}�g_�|�� �̸$�<��*Pbo3`�Ĩ���|�l�����?�Mp-���-Sͽcۗ�o�a�Y2��j�͇���/O������	 �ei(��D:?�H�$��M��Z4\�R[i6�f�b�){-O/�����O5w>�z���G�}P^��l�ޑ#U��dNx8�|u���傤&��3����rfQ���2�c=�b�.v�-���{:�֍� Q���L�����dǲy:Q�AD����|�+�&�b�Dd���Hc��GN��dE�����XE%���O��6o��!�A���-^�U��:&V�K��n5n�2�_��z+Bb�J[;�,bnf ���.�_�øZgR��S����G�XgG;!/_?TG�%�e��$����?��5��N�
�ҥ���A�r��b{�2� -%�P�3����y�T	�3�kǽ�<6JE���r.R�䅇��P QQV\]R*�n�y������P�"U�]R�C�}Z�J����jڱl���d�H��(T"�a'�w,������[����K��0����NI@j<��R�Qp~.ۦ�rI:��7���"��z	BV����)g����8���}�>���/H�k��������� D�^s�1]�7���{���Å|*���k���@`g�f�%�=)ܞQs�fr���l5~'���$�P�p�!����~�~Βtjp�b���Y�N�s�2�m�g���O3�5(W�1x������C�j�q2	��F�����2r�sY��ؖ>a�5��`_m�}�!�>������\M��8���0�2�ׁ�릑�]ldn������ap:���t�P$h�Ap�C�a�"Q��>N�!-�V`
�;{v;M���VF�d���C���^ǐ�A���0�񇒸�zjtj��qU����`uQ��Lनb�?ܺt�xa1�/5�_#�F�s��J�I��A��ߧͶڀ�y1^� ���H7�G�C��G���yt��l�QA^m�����f'��W���6O!�7j��kX�PP�XqNn��'Q;��b/���|&n&���Ғ&v�|�}��n�3���^j�鹐�k �k^f(�2��	V�q{"]?6�?Zꂲx��x���pMoLm�Ri1��'Q�t�ЖPQJ#�
�E
$A��8�2�2��Oy�2�z#��v�:�*��b�2sWW�<��dťo�1�k�;H7s2W�����$�P�ȿR��z��ʬf��1�N�d�@�{H�� !���h���[[)��w�ӓ��g�4'�����^L�U3��.������B3�:�YW����{�J �vYyG
y����E@���&�uMu�LW�|F۩��¶����S�M��_�;̥�G������|qT�"!<S�b����l�����W: ��2[��L�]@�h+����ڃUst�b'��G��.���g���
b��Y�&�0o��'N{��A�Z�t��J�Zu��d��:NR1t�_x9�8m�4�Y��:Y+�#f�����b�b�\�+�n�ͤ�bWu&�ן=4�B9&ğ���ྑ1��@G�H5S�����
�ۓb%o�A�;`쉽���cwvj`�$�
ʮ���+��t�ޱï�k�/
<����k�D������{�h�>\���B&�x�[e��%pv#?1�$���#�Qo�QW�~���"O��,�_���Օq ���B ՛����� ���dtJ�~Hxķ��0������KbaV-�g��W�!$PI���G=��w�~�2'�,����(6
���\ݻ�d.��z�_7Pd�M�g���p��$�a�_c���|��(��U���g�z����������
'��8�ԈX�B^8X�MW�,�:�?7x4�o����8�t�s�s��f���W��j���ɿ��
��?hg=1�'@c:#�P@���z�ཌྷ[&�� �:�獄vHh�u_qH�1_���F��Đ��&��Xu�T'�Bt�53LfT�ɨ:4�+�p^^��^́Ћ���K.���t*f�n�z_]�|�ɤ��D�O�*����W�<����%�z>\h՜�{[��ml@��B���/0���p�;�Md8��oK�|W�&o�G1FU؜��rH���6�|T�VP�G�[�+����S&���7�ep�ʖG�yMT뮊���J�h�hv�/+ ��܀i\aO��<b���#��B1X=��c�z}�|�W$�Exl������l�#�x83�h���!�YߧiT]u:إ�t㗌��/B]j���w�XAقTp�*�RY0�)}��K�5���B��҅$�<�t����)xV=B$zPa(�n�5�
�ŤX{f��\�(�T���]a�l.�]@�����᷍��J���k�%�E����!�vg��@�H���a�TlJ�[�}�]�S�g\\��GVaQǾ��r����-��Q�Q&��'�)�D}��Q�q��v����fr�o��8��5a,�(�/}Y0��剤�ɲ��bV������#��k-��l�������E�H �^�mO܆0�H��	�ƭ~8������p�l���/k�G��l����In�}J��Y�F��Za�  ��K]㻝M|�K�'z6��yx�!���λ^�5��И�>�S/��]�vvr��u_0�X@��J�D��%ff]�Nbm�����:k[=����a0�H-��	�ξ�fN��U/{n�^�h����Lw�HT�|7t|�x�?���'�\��Kq!i0��_��NK������9o!�q���t{�L��1�1�p0�O�N=��]���8� 
x3/�,C'�R�:%)H�_��v8w��\���|�����Rl�,��%WW<���V��ci�Cu�����!���r �Fϯ�N�;�y�DL^ s��i����T��?)z|����zbs8!�ޥ\�u����+�žD�;���e.6S&h!䒚�"D=,S}ދ��.���e�E 4.hـ�N�4lw=�P\<�#}����+���CF�K�Ru���g�~���)�ad�D'�ˮz�-L<��u<?N�rP���1����+Q�+��s��N��@��25<�� ")o\�HL�m��pӺvrz��/$})�r��qH.��9�x]G�vF�!��c>�1r��R�NE���	�#9��Í�$TQ�K�
�:V�q=M˂��F\Ӑp���M$�$9�f�����=�Nv��7
����p]��Id�x�Q���qI�g86S�85�>Y$}�L��X-�'�}i���E�
@��~ހL��Ɠ~���=YH��7,� �R���"�,�lt�`��n ����b��J ��.G��-�,X��Al��v
�QA�O,�#Z�\�(S��8��j ��g��u�����@S*	�0VV�`q�p��l�D��b���iH��x#r�\�/,��{t	d�0g�hȧ��]b1+0�k<�_�_���8��'�Kb��P�_Y5'enW��pE�B5L��C�;���Rĕ�{�`�3��F����Ei��]T���Po=W�"�/⑳��V>1�#�G��o�~\P��/�RjZ�!��o����\M�"�����G+�@�?R���4�%�KqӨ.��Bk���N� xc�q�RR�^�s~�.��u�~��t+�/���ĶJe<�@v�<D��])�b� �0�S�7�yWJ��򙮻㥑��8[>y@��[_ú�-S8|ǖ���خI�� �fV�@��
������O����/����*�L�Nn������gH�bɁ:�ߟG�|-wu@ǀ�wh��Z�oN�Q7e�Ⱦ�z�|q`��uJ�C*�M���z����@O����'�t��7�O�/��̷�~����ö���s�I&����m>v�z�i۝M�0d�P_I|����1���db�j����qb��ی��,��|V�h��W;E-�r�G�z�'7q@gZx�]��_��:B�+[Q��cq�}}P%h��#|�;��]�(|��a���[�o���>�g��Z7|�yq(��$ԦY���I�ӵJ?x�Md��4@❸��tv;@>��:��,��dgR9�f�ذ&2nd�|��mNTF�
~Dr�v�iD@���< s@�XM���%��)�\��`�����Y�G�����̢ۿ_t��AE�~����d�y��l%��R�~֦*SB�s��Ԯt��͝yp���*���!��SV
Z��)����;�l��,I���2����/��s�L?mi"����'c:�^| ��n�|��I��&�q �r�3�G��=đ�o��Ϝ9��cF�5���'�L��䦺��xZz�<}^�;�3"tD�� 3�ͧx���ٳ�`_�/�w�[�R��i�E�D�8�j�`4�s��_�S2��X�x"M�%�S�e*x�6٨��<"t����p�G�Sacc�X�n:Tj'�� b56�	��v;E�I����g-�6-FR�N�ꯋ�<�J��Q]��3�3�`5꧝U������-y#Z���D֙�3�Zs��᢯��%ؠ�߸\� 06�p!�v A��.�Ө��%��'�܍��hݗR�89��˃��W�bF�`?����S����3���d)`@(Ȩ���F��I�}	rcdLޫd��=e	J��B5$��@v�q8]ec*�L����1�&�r����/�Jp�XE� *�"ͫ��s�a��*�eq�����x�L�\؝�J����P�a���3},ث���k�t�l��d�:G�%���~X5
�˃��£��!bx�ַ?V�r~�T��wʁ��E�0��rE=��Zʷ�k���]�)���l�jV�R�M�t]�G�>�u��6`ǁ�D�~���g�n�J�*�/+YV�i�;�C�DX�4ҍ
�\����Ի��TJ�������"�/�=�s!*�o����-	 `e��gN)��o
�k#�� 
��V��d|��+k���P��{Gdɔ˦tH���t�#��C%?�:`)=�7����X�I��X=�E���tsZ��w�N��ϢV��+%�����H�}.��9V%���L/�#�E�݇1!��������b�:}�Y0~mf�w(�0x���E���|�?X����"��\�B���g�iN�Ց
�Bm>�������ZV7E�r����4��酎5��{L3�|q���J����*&��MS�������K�E$���Dm���y����sSsz���HH����	���e�|�>d�ο-����{s����T�و��
'\�K��d��+F�F.n�\V��/��
 ��d�E1��rj�u� �p>C�ʙB��3說y�ε檼�'#�姴{S����z �d��f̝q^J��f���8��˝�b��@U��_jL��_�hKUe�˥t�M/\�h�qu��pO0�>��SD��LO�x*aU5�&��?��Dl�S���C�+�_���%��\Ȕ"��>�M��ٲ�ՅXO�>�-���]��B�yP�)�|?�[�R�P��̈́4��Ar��kI�;\�M�۟���[��*/.��U����^�(�Z����8���(&l n0���}�l�>�Ւ�}�Ӯ�EWi�Z�h	w�b\��i���aZF7�/a$Lk��:��uB<̊�M��*Ze�@��8��Pv����c�졧l1L���X">w2@��"���������jU�~��p5�s�	]n� C�`��&�z��M̩�0�j^k�������-/�Ur͜}Q�r�ܑe��Ą�BP7'逇�<Y�AG�H�N�(�*�o��P�}��	8!<�pw�B��I�U
]�c@���w��u ZWxGJ����W7� ?����ܧ1��ջ�'=y�� h"�¹�~A*��
��y �4�O�a�Ȝ,�H	[�}��F�������3s������j�X̯T�W&9�׸�Z���yD��\H���<b{��T���E�צ��0��袘�s�����b��G�^-������Z��"�RN�_�+��\��ص	��4�O����LlUݼ|KY)��.�Y�9y�]��`|�F���p_-�Dl����D vfa�@ᄻg�����P���}]Ĳ�	$���f@�4�`�&N��,�R%%��>r"T���;��F�Q0���ㇾ�CݣUD���0`T���߈�H��2�q��TO7�=+y���ލ�bO�Jx�K<{����Dx-U�a2v����,�8:��+��z�P�G&q�S!���X�bB�Rڄ0	%��������aa��SL�i�*��2N�9?0�ˣ׃�Sߥwr|�x��� �5r ��ϟ?��	���_�Ə��݅\����w_���<�۠���5��i��}�H�/ѸA�U�,���������h��Ab$b�M|��QV]�0�rځ�m����q��5:e��n�}�nk�k ̢�u_����<��}���a���ДH��[<��n,^K�X 0<�9J[7������ 9<�<����yM\z��f i#^v�s�}��<`(M�������Y�������@�qV�4��[�C?��5�S�����u<���gR�	������Pj����	�(su���Nd��Ƈt���K��<��h�8��ކ��`�7�9'F+���Yԟ� 0w��1�Yt���^��5o�G���v�F��ʽ�����%������=�]|���FY��۱��6�����K��Q�cI��N�h�3.5���6M��@J�̓+�zA��:kWWҷ�*��?�����b��:�|�Pԛʽ@r��Yeq4��ǈ���M؇-8+{X^H����溆&,��yT�����pg2���� ~��)�k�e:�'v S�y���П�R!{���R$xe����t+�/l�ݷm��,���I�
e\��d K�^��TP�צڹ��o:�y��"�v��˜,�Y�;�ON�;��Zr��}���.���9���9�t���㉋ޭ��Ԟ�g�$�]�P�>��&�ߣ�0��I@ !���)H��R"�֮���iq1B�ܳ e-���ï��Xֱ�_�2�T�IV}���	�r�`H5j�ory� ��i�<�Vt����>���|��h6��z�&s��Z�b���v(lV�c�x���D�o��^�QsO����E	���2�5-!�\�������yN8��W���m�ڴ3�usp�ʎK��b�?^i݉��]��k���{�)�l�Dɡ�㚫�ԗq$������%����!�FZ�>�g��k��O�.JP�J]s�|���o���T?�ʻ�AC�Q����j���-�^Z�A���d�#O���0�h	=gQ�y։>H^3��O��Wj,���
��.{����M�$}TW]9/�^��t�' �@�ð_E�@&S�+�?��~�~�H��H�2:%�=E��e?+x6�q�w~��j�w�^1f��g1
~߽0��4u�'�wJr�Tŋ��-��?l�at|���թ��X�JPJ�8bjj"O0j�.���b��į���#f�-���{����XH ?+H>/O!AW�U�+���*�8H�c��C�!@=�(&���X0�A�8Z����EJ/6����kK�!<#,��l�*��R+w2?�ki%��;=�6I����JU�"XO�,��]�|��P��`��d-NZ� �P�}q.��1��^��.�j�Y��Z�Z��l�#��J\����A1
G� ����F�@����=$d�_2fq��s �P��=���G�hC�$+���vc��
�W�J�߬�z'�г����(s�ɘX�5�%�-_V�&�Rb9��F[Q;<z���Fkݑ��X��h��]�F��y�g���x��ږ'�2��c1|I��57���J+�޶�`E�#u�n�k �)�?�A���=��?y��;o���̡���Z��N	!��=��B�k:[�K�ӎ
!$z�N��y+"�j���lQ��b��/?3)�lK��%0�Ū!�x0A�Da���	��io���
,�G�G`��/��.�]�B<�����!׸�M�W����������-���ʟ =�2t�x��∁��M�X������� �g5-w���W5��HZ�lh���u(`����Y?��+:PC�D��ꡫ[+�Z'F��A:�N�'6��9�/Y(�"����;ܢ\�����:P�k�i�2l��Y=Ib�S��
��9�Fv�3';�
�߶)^Q&��,�]�..Ͻ�Q�(K6��.�A)�N��*e���Թ��K#���W��1�ø����Zm�a�I���=�b}�	�������L°��] �h��J�./��a�̱-B�]�C���bC�(�?Śxp��gCk4�< =H���1Z�.~���juQ�*��d���E�ח���S��|�n]��Hy0�6x���۞ˢ�b���(>j�v�+��
�����~��k-����w�_s$�����F:��8��5�ڏW�����Z����pT�Y�^'������&�0/=@�b����lrg~iD�.�C��i��n�63�_���Q���15mi�%�T�b! *:���n 	�Y����lpK��zqW��d����wQ(rR����YJ�`�A�ެ���b6{ů3=.�'�Y�r��f�1�:U�[��VK/>5a�*�0�3��C%L������*�
����I�������2!w��~���|$2���(�	� rm���s�� ��gp�#�Be�;Ѯ+lΓ@���3J%���;�%X`19<c\����Ipz�,�^�#[LC*��(�@����ʁ�8�>j��Q�,��������Ed}?&_�>-@p�q뙅��E8�9j�:�OWW� U��M��Є���u�U�w��wL�\�f��I?���2��q����?џ?��H{;���������eaocsAb�^8Չ=�0~�nm�sm��|{.�Yn{�ўkA�`9��#nҋ��e��h�W\"�㻱̑v���R(��Z*c���M����0����aT7s����>�?-��_�8�Z"�ȟ'܍��:���.G�RT��U���]h�����/W�/��%�i"�w ��q���B~ ��uY"�ۘ �h�.�,T=ʇD��p��@tG�2g��oμ��� T����fv��ن���+�n�ӽ@ɃE��4�G�(�M�zV�U�'gKֶZ��%c܎ET��[�xux��P^"M��@�Ǽ���<~��1�)h��D��m�(�y�8��n�U�����^�3 �*+dHW	�Vج������-��9�<�[��'�5Cl���x���6cN,_���}�!���OI�ܬ�M�MpO�����=7e/[�]�#!�?83!��5	�vM��w7���ˉU���u;��0z���P���k���2�p�6r
�~���u|A��-sՄjǮ�R���7�~A�'�?5z�@R���;� s���2"c�#-�p��Q�&���&v��'&��Hהe8�2�"c���Cf�z�.�4y���U��Z�����?{�*g�g�P�aR0iH��nrj b��^�Ő���*��<�hfNp!ܣǿ��xY�SuXK�ў�X�Ҙ���,��.<������r����kV|�n���dk��5� �G�f�	>�)��t>ԝ�Z��y�|�.`a�9�'��5\�DK�&�&S~�� yn��Q�
�0��#y�	rp%Pڭ��<��]�&��p����	�jjcR��y���	r���w�d��'-g���"�|����*ޚ�+���&r��4�~����}�
k*{�8��}��[�.4��W�y���`B���s��D<�[l+*�C=����	��}􏾶e�U*��u؛d��X<)��\����x���DK���}w���%�A�5���)���=�=^�u��0�俳��v�U�4>���ע��xa�&D%QP	~�vΆG3�D_��٣����(ƵC��cۯ@FE�s�芄t���@���M�ʁ���Գo���w�=>/
xpvv�[:�+�����2k���>˛�;�@P e��D�J#(��=�FA!	�
�Y����nnY�t}[�5A�~t�2]U,?ٮ3�P\����ۜ"5���#����y�k��0�AE���� �4;Qb�x����{�j�����z4R�}�`g��
��Q!®E�E)@u�
��p�s��KI$��q?�����hD5�p,�?T$��o�:��\��B\종ɧ<��;�����Z��o�-҉�w�^Uǻ�&��c{��Ћ2��+j�=���y=>0���!��kr��s�)�wU~.�a�p�E���V�-i�oHZU�D,n;��+���K�����c���k�q���[k$�c)�{�rbj�C��@�\�l��D���5(��/��8��yA�vQ�Gx\����s�]g8b�@Mx�����!�@]�z�\!�t$ę�u4���Q��(U��v\<� ���M�8卾 Ԇ��2O� j�cbN���hJ�ͮ�T��6���^B^'����󸽹.l�GU�y�n5 �qa&O�K\ԛJu�����g�DVkq�B9�"�]�gz@��_ڐ��=����>r%r�Ut��1�N�G�z�������U�O�=:I��tʙ��� uݮ�v�Hq[<�}`��í�g�)Wv�|��Hk\M�K�h�|x�$��\�x�����a�UO�2�������L������B�c3�n1]�Wt��x2�{B�g$d���1�c?0A�Y(�1e�'K
��hm4C�r�"a�üN�!�`�9�W��0��N�\Z\�/��P8�P�� 7Ys]�8��y
�C�p��r�2Wdkh��"o�m���A��_5~R��W+b����=�&���䫟���nv��]܀�<D�����6޹��v��9D��I�7�Qv�,�@a"X�j������8-S�U#�y���6��ޟz�f�4���$�]��ܿ��P�t�a/ ��d�Z�jɔ�,9�>�|3w.�g?s��dT��"욄��'��jڅ���ͺh��e�+�P��F����;��=A^��p�I�n��h�,���1����Um��4�(
�B�ܚ��gC]�.(�~'�r���;��I����dB��H�׵�1�.h%:�%V /������K>�������v�K�ǜHNV�0��$=RFgo��Ӌ'|/�wC�\��r�Mp|1�1�`�=�L�:PX�\�1�	R&.Zqݤ�����J�E$!���$��9b_o��g�.�QT�����S��A})�&�km&걒��ٲ�ҤyG�tn�g��V�WS���A>�3�>x��X+�++{��d?��+�4{�Mփ^&�X߫Tn�hL�Ӽ�M#�(�#L�w�ֻj�p���6� ��N�u�4����4�j$�+qS䒴�GN���1�{q0R��&N^��=A�H.�L���>q���I'��Q�'\2�.s�}�h��E�C��'!�X]�u�����ʳ-)��S�4��y:��j��z�S������}��o�.����Ђ�����##'�s�
��\�\���^��E���д�B��_Y�{�� >�1#�A7E��Բ�u�y�	��o����;���bP�q*$Z�Vr�sYF�b������Ӏ���
&hM�O���8�$=S�ުv�$�����g����l���bT��;F�osUg ��	�3��!c��zp��F:��ڒ��*��bu��bT7�O�_�����:�l�/H��
���DU*��OG���� �1��xf���_����R/ ,�qg�D��|D��B�U�x�k.��s$�tN� ���8$���]X���!�r�?w�f�$�e�2\�I����p�a�L�����''::mβ�}���P(� ��ė�,��}��� u��p��D�W�duB"�p����rќF㑉�<y:����^���֐-�l�3���bpìX�Q��9���
���&A]���-j9*�S��;�DHl��� {��<��O��rb���m��'~�(�(��fX�qG�P�d(�ն���s�zl��l��b��|������1k�LSW�3͓l�в��_��i��`�V_��l<�
�O(���G˫�y�����څ׺�4P��u2�+���5�
��.�(�8�}�R���B���wX/���!���Q�`͜*����/;�!JP�����L/��z�/�|xtU�vi:X�A}Q�B�g{��=,2��L��ER���p�2��'�|��V�(ņ�mD���>�KU��Ӝ� �cqOJV�)m�?�B�a���BD$� &^�e��-�5_/N|�������E���&���h6��4��C�rX�=���b<ۿ{��mSD�*U�
=Y;�����^�W:�� dZ�1��)����`UH���ߥ.my6��'k�z@s����$Xq��%7�<yQ���6;MH��h�L��*���o�,����>�2��zt>�ɯ�a�8�>�a��&�
��ym����ߟ�z8�L<#�m�H�!�"���<�%��{=����0h��O�"એ�)��C0��C����I�܀�hmL�������E%R�@*b�h�i�[[��RtgH������nR��ś;� �k�V=����"���A�RqJD]�R��heZ���dcbW�?���Y�R̩w�͋�':���M�u�QbV��z��`3�p�CTm9H��SX�?'��<�D�L��ٴ�` �U�E�P�q�ISq�|�KQG�����X��P�g�K�g�M���>X�qԼ���A�ENd0���s�-A$\��2��ϗkf�|��l�9�^<�*��k�Jm���>�k��Yܷ���LCD0=t�����6��_�)C�>� f$��B��'1�5���.�X��J굼�!64v����frn��n�*!���������[�7�M��}%�K��T�4�E�8�+I���U��a����.��Q�׿���X���n��@�������Aɉ���gu������){����7n�2x6\_u����Q���32��k�JM�lp�������n���J���a=,8n$������o3�BC���^�\�6��e���&Z�3��%A�*��Ѯ�*{�
)��C5$�n4|��d�����@ުW*�O	^+ĩH�����n<���n��`gM�����_�Cb�=9�䎠#b5��'��k�-8��)7+�۸�0�=	d��-�����8�+9�	$�n���F�#�!|���i�@c"m�l�Bk��F���(7�/Df��"�L�n1�:G(�RT����:KN�2���C�(��Ue�ZT$T<C�r�X+
ȯEY��E�1�u�p�nTŵT���1�,g����k_�6$��2����Y�Sb�@p�Ş�����h��:�ty��~gI�u�&��?`B������h<�q��H�n�#_�p�-ƝJ,N\��=o�tn�5����0�p�K�>J_[���L�Ņ�O4Df�� �6���N3��#����9Y'>a7�^���vf�8��>K����m�Bߢ]�Q�sɥ�f7�r��#w���.^�� u?�\~#n$x,p#f�E�
��eY���Wf��q����7��~bFrG�����w0�:��96~�xE���Z�O�EYr���I�����O�&�6�ŷI��P!"�6vcS���Q�Ph=N�~[�H8��
O��gi��g�fg���D��ӝdeϰ��v�g��CkM��j����L�tN[O��O�a6��+S_%ﺟ??��p����g���qt��Us.}�����j,P����A���w�uew�1C�"���^
�����*X�e��A�B��'���#�nJX�^;�b��i����Wl����Zo��2�}��^���2O�3��U���1�EC�E�S~�&�r~���t@��������#�־�i9]��1qD�.���F�oR2\l�������=�5C[����������f��zq��Op��uI+���~�,RVB� ��F��0Y�$�`D�}�mi�J��u��@��+�\��H��/e֔V�i���3%%����-�W�жh`2:;?F5l��B�m6����`I�����62;��e�O�G��!_ONV!P	��g�VprL���R)N��=�������+�=�%(J�)n��%�L��U\N�D��#V��\un�2�*��޾'0c߇��u�H�	>Ӟ*��"T,y��㗪��.r��g����Ղ�9���x��Ō�O��嘆c�}h<תJ�l'7�l�={����T�<9����ł� a����(����7=�,��Y����i�Z����s�~ð��:��3@�k�%do��wͬ,��zBV(�fr��.^�	-Uk/~
/��Q��T}��d��&��1!�_�� �w6��?+���BaC�RA�����m��J�E0k��s׭c~��9{5�7���3���Pɇ�cA�҇�oǉ�L��f�B��� ��io���n%�U-t�G�q4(���,��L��T+n��9�W��ֶn��З�7�����9R�B�{�^e�pK��ީm%?�N��e�6�g�R�0��E�
� �I��]ً�N�w���kڍ~^=��%�Z�����������J�П_[��2g��R�غ��j*Q۟J��Ӎ�в�������~�4���\�k����޿����&����Ą5����Q�`�A^\j�}E��ɟ��g���6Y�?!��iu�.ɴ����[m���e��S/	g���88��)�?���ߏ��A�	�x~�ݔ������4��EglQ��O�5����9=��+��f�<'�b�:�t�躀h��R2X�>X������k�I�6q��v$p]Rv`x�O0E�x�wX�٩��o�"�ު��D�c�F�����0�� �01��^�ȴM��gC�9��h=�ڼ����K
�O��q��
_��q���W�Z���\:��ѝ�Er���r%��c������ŗ�Pc`�H��,��l����i=�¾�pz�m�Z�m}�$�Hrye�:8�9S-%��-�1��<�7���z$&'�Yj��ݞ�9�%�(!�I���:�SI��uw�c����7�X}�K��N���dLŴC�?����(l��T1+O�L�� H ���(6B�I�ˎ kv#���HiGMw@��q�C��mCJ[���"g\���|�B��Cƿ�Oă�5Cc����R�?�Y�c��}�MWTt�k!��zT��1�.@ղ���{$^�S���`��_p��Ñ(��k���I1[nT	�5���:��V��m�l���ש���A��}_qH����ƽ\�=/�����Cr�s�	�E�=Nq���؀�ޥj�-�6[]�t]�5����M)��ܸ@_H-n�B���?�� |����͘�=�fY�*g�gac����H��� ��f4�����^���\WP>B�,�:�cK� �L@L\�bB��s�E)'T�����{��e�_[9:�}~{\} �ؠLo��������^��AD;
�v�n��Mf�=z�84�n	
h�Cy�+tu�W,�_\�FP�������O��������#�}$������%+'���˔��B��B�z�ns�Ǻ|8���r>#�ѻ���}������p'j-l<����ս���EJ�(lz�7I��B�}�'SgR�k0S@�W��M����]�ܽ��:�큫P�dw�'�MN�N;��J��YخHTϑ}�c��`+��B!L�e����`Q#ˬx�ZP��)/��,�E��V��W�
�Ԭ�=��E׵�	�G��wV��;�6{���E���M<��nak��)�`K���w����� 4�]������۳���^��"d�/�S�=�4��btX� ��C���쪳�,�a���!�'��с�m�-��(N��Z�e��~]SQB�Pl*9� �x>��#��n�>'���3�h�j���T��#��c�o��Y��vv�B���1U�ǁ�9�{�[� ��}�e��Z�p7��<(*TLj$���[�#���lA�ޱ�q��`��������Sf��K/�nV�9\�7{���HM0{-��b�a�#�� ����%9/�\0��hO8s'��3��(��K#zh�=H�����o�I�M�A�f�KnX�ЬXW�Q�4i"R�O���?��q�f�[Iva�S��,]je9�h)���9��	�`T"�I2�ƅ	X뮘h�_賨lH�9�́��i�h���e{d^|�ص�q_0L!:�&y<��d)�,]��,���h|�T�{�OZ-�"ѢC�ʪ�������d�f�O�s��]��.�&$d-v�]�	`o6%�l�;����2�:��@�7����	l�vu.ltq��5�,�xl>�Wz'�f9�,�����¯���^/��*�T�c�\"Q�]o�_�����9�0���%nߟ�z���)����nO��8��2o ���GXa1>Ѩ��⨏��=C� <"b*�\��2���ȕ���ZI�ۘ2��p��)P��ꗹ�
E-�g� ��h)�*�c7(���t*K"J��R�O��1�j�1�v�n�m���M�G��q�����.�ÕI����k�;���'���&=�����U,*ע�
7�~�_��Mq�}�=n9����ۥ��c����_��ӌ�P⿦���#%5��ھ�E������޻����E��/ql����:���@���q�?rAg�U,���*��;lt�8������IJ�>�u�'�����2wG�2���/���5Fk	r�4N�;B�L%�6��#Ά�������9Q�i1�dz�l�-�˗��w�� St4���������z�^=���e�]9��W��Tk?ox���7ZO����vID�'.���X�3�j?#	��cJ�\v�#��E!O�)�c��:�K" ��e�"E͛lr�B�j� �w.j>��SL�-Ѭю���(�Aɬ>b����#X^�p1Ą}M5o���jm��L�a�Pε3I�*c1�1���N�����m��8RJ��p�~re��o5�3��/d*�9Ґ��n�R<��m��r�b���<�v�k�aV��eT7��5Y�ܶ5K!���K�te�jo��B?d�w��b�p�����
��,�yUs`�K-���6��Lo�S'�B��VH�ZQ�p��_eͬ��w�k[�m���z~�8�p���O�I$�s���O��B�fέ���mlL�)��d��ą]�j�'��n���K:Q�XjNeգ�6D+��ڵ?6�g�j��ς�h-�7�kԆ�g����v��z��G���[���#~�|�e�V"Q$ڪ*%S8�e�l�+�2tU~X�g����[h�#n�&���~���!�m��s؁Iv����L+�Hg��SK�`������������>��W��s!jX}���:$�s�9X��0��*o�Sx��Y�l�:�C�-Rl�ߗ^".��]��u���8f,�n�}Z ڊf!�am���9M�7v����ԃ�~ۚ�n�stf��� ܻ�9�j�e���� A��u	���[^�NB9T����v�\:\LH>��ܘ�ۦd���I��|9K-�լ�}��������/��S:��âc���FӀj��!<�U��b^G5	�4.sˬ9Z�D��u>T��͒\�ϵymL5�9���7��"��NX�aF��[����#p����L��UP)��\��[���h��?� ���_��F�ZrX��w��3�>ń�2�/�L�hv~_N2�C&��_�����`�Y9�Jw��h􄑲�s�@c+�#����D����ѧ�G$���)X��LXd��m^��UD@.�������M���}���I/�����6�d���/����C׭���
�НAA�<��/
v�P��h�@0�@q�d�"�(����b�5Ҝ�~c�k��g98��#^f�Xu�� �rʢ��A�'r!}0��O�~H��d�����0�����>l:?e[k�� ���lS�]�����"1�g� ����W%������'����1vHV_z'��6v�$ޤ�ZO_�Bf�tҊ�;�k7��ʗ���!�TC���C�P��ܶ���,�h��(�u�2	͜x{e�3J���k�[��j5T�Zq�\(�nI��,����✫פ0��W��+�/x�F㮨}��I]�TJ���[Ѷ�K�"q#�`���?w���U�g�!1L��K����-�C-".1���iی!���Cͅu吶~����[m�YZ;J����V9����&��e�&�R�[M8�H��ړѕ��<!C*�vlȂ�D��։�����uT�{���/��W�%�'&���|5xgOXG��2D���d�u1��XƠ���Ll�@��L,�*j�^�X�ͳ��'�	�K;i�����X���؋�U�;�,�Չ��߶�e#UZ"�jn��;�%�g�(�<�w�hl��&D���c@7F�	�Z����{��}<��7�Q��c7�ǎ+ϊ�'���_,^b"-e�jM;_&mpl�n�`�`��6y')���S���?���E�(<��j�ɤ�b]{W����λ�R�z�~�	��M
�H�Z:~TjSv+ݡ��~&?߲�0��tD2�d�[�{�ɻ�j���~j�h��ޜ&�g;�I+�Z�z�lL^
�۸4�:���|��鋰��&c]�k�"��N#4��Q�Ï�Q�KFd�|v��N��\'�� �px�u�������O�{hӉ��5	����G+��Ƭ.s�0m�_�R?#�+�E��h���xB\G�g�|�~"4'�H��,��~�¢�M���E��}M�����#�2����A����2�"��&/?N����g�H.���gRdww�b��ǀ�Q�c,iE�-X��m`er��8��"����|.щ"}��C@O������zV�"����>���⢌�@�ܢ��n��5�6O�R�C�'i��>�|�b�-��Cǃ;W.E" �B{B	eD��	�g@^�'���O.��a&=�w(�*I��6M�$�q�Q��9uz�����9��	�gW�~��}JL�!�g��;��	�v��.��:��Y��SG��PC8ˮ20c �7�ZGP5_x�ur���C!������������,|&G�����p$�b&wf_�n�Q�Hd�K5�9iW�|��ja��j(+~��'�����i)��:��
���D��C@)����!�v�r:�2jf���y����W�Ȩ�Ǣ��]��D38����>$渽ӊ����f������G�����L:��y�m_
�÷>0�������K��	���0]>���aԇ�ya��*�]���	���t�L#�����y&vßQ�����kE�К7�J>{Qu�z�n��Ͽ��~����~#fE�)J���g�*���M@�l���{���%��;�aJ�C$i����`(�~?&/ag����I�Ɯ�ų�oL���Jd�:L�u�
�K'����d>]Z��ke'����h���	
T�B]��F�ÏY��WF��R5�;��B6���Ȗc��I�т8��NQ�e#����]%�o�X���A�������=?B?0:����B�g�Ou���>���5�ĭ�p������w��U]IM�s�V<��(c�'�����K�7� ����M>]Rp�M�Tv��v�y��[5����Ju�YyF8$�]~��b=�ґ����I�� Th`H���q~�8��&�iI�:�b>����n��G�5�cE@u�L����zH;Pʼڕ��D�(8���!�#?0�,�֍���:M �{�����&�'��f�v�
�iCҦ#L.����\]�T�AO���p5u�^��Ԡ�բ��t<?��o���KP4�
�P�K1Hz�M��Kf�
���G���u��X�=l����}G��=�*����� �x�.w�V@U�iS��BĤܽ�C#��o�D:����1��qR���J�ޮ�m�r��A�Iݱ>x
����X������6��@��'kXu(�����I���������{�y<I��Q|����h5��J>�l:��S����c�Nңvza��[�|a3�@��_����b�9{X[�b�K=�TO�4y�)��o!�TCp����g�5G�H;�*R^�g�%л�1��	��77T�d1�=¬Y�	!3�ۚ�p�T����G�l�ۗ��g�1��Jg�o>ŷ��0�&��3�����"���V]+��j���f�^>�Z��P��,��?�Cq
X#ѫ:/�r �Gy��������`���>F�Ƞn U���!mV٘�8�:l�S3�2+?�A�w�]�����s�$5&�̇I�VZ��f��4��?����b�XNs.�A�W��9�ݑ{�|�f�k=ey,�v��(��=�W���k�R�Q��!����Tl�;� �L@�X	��8čB!f��k�;򋗼bT�?J�\Oy�f��ɶ4���Iv��kP��# F��::�����O��+��tvpp�<��c���M�d��]l?!-�Fe�$$n���J;�����	�)<�%2hy�	�iͩ���6d������}B���/۵j��?M��*'����&�bĹ�HȘ�����u!HʳR�Q�r�=���.'��Xo¬�
2�%܋�Wd�@�s�n�4�r����Pq�$gQN�	��K絕R�q�S�^�(h�.��U�;��������� ��P>���/������t\r�w��j@�V��Gmx�,�$�O������{G�aBL�[V�6[�xI%';�g�PtX'�O�Y.O��;�)l#�H���!�K]� ��%���:.��Gi~�3[P�ک�`A�Eec���>|��B�%�&�A�52�����ݵE{�TΝ�KZÅ[HO��d���;�������e�>�تn_�Z��:����P�_SóQJ*锩�����ߎ�4��Щ�1�ǕȮ��H��`�z Wu9��?�V�������|���C�]�~���9ح�j�&ֆȨ���;)� �5u�G����G�&�gM���P�|ܴ5��IR��h�+�[vc�-�ϔ��/n��5Ի�.u��n�f���n��h�ڷ���Ba���u	���ڸ�kc3�V@w�Tl�Ҡ�2=��}*��~���NV�_�QY�4��-�?�v��s��^Ӄv�z;��z;��қi�$�@�ld��.������#ݍ�m�m�?�H&k�*G��1݅4�w����ѫy�f^^��p�0REL/�m5��i >�\R���Nۃ���Q��~
��
04:H΋��*��Z�4:{��{�G�;�[�Po�b`2����˥��sJ�]*��nY���`;`r{/��2#����k.GLI�?]KP ������̊",�^G���>��J��M��z��A
g��|&�W�Y!z�H����"�2Jt�}�&��4�3m5�5�CA]���<��V;����@��Ra'h�.�f��,�*5�3KQ����t����_*�����𫖙d唄!����}���'f8�4��x�S��"��>g"hk|M�0#�$W@VT�Pf��^6�H� ,�WA�,LǕM63�X��	gI���_�[��+U��T�M㮒gF|�0�������4/F���^}�R"~��.P
�k��NWx�$��Xs�x�r��u�;���AR>+y&IY� p��Z'ʭFi�7��Z_f�Cs<�E`:wp�f�MoM�Zۿ^W'㣟�"�S\N}�]�S�:�5�&ң��W�=i�L�z ����DBf3��ӞfN9D'�ЗwT@5����j�V���+�Aʢ�-6|��g�M�#�W��2E�9��fA���
�r�Kßۈu��	e�Iv��25:j�6���8�8���o��V6�B�6���l�{@���X�@��
�z���*�N�@�pX`�]8�6k�0����Zx�6�K	��W�1� ��|��3;O�v�
]��Why��Ә��P_��:�+f{��?����y�:{�����x����1�j����%t�Ag�F-l@�tV_�b�Aַ���y���6��uƪ��⌯��|�����&L��Vi5��g ]<�i�W, G�2,�i�k�"�|9�پyL�M+�n6�!���!�B,�Db۴��tj�򶅱.|��r��:_z�Մ��&�6J`*��:x��P~kxV�{%�q6�7��8�b%"���"���v��$1n����F��j+�`�mq���Q�(U��v_���_����1�јQ.�
���H���&Ć��������'�#�Gy在�*#�
`�?]��p�sʛҜ�$M��������e��X��?6HqRj@pV�j�/7��y���]w�j �:�K��&p����.y�塇y���'T��FI�,MM��D1$I���MW�l{�������TY~c�l�ޒ�h����{z��0�� Ͷ�"ej� ���'���BG0��HV�B�Y��W���f4,��]j�ĴZ��b��|U�3�z�m�D��V�4����ɱ��H�����E�B����3Y���(�*��>�9���xl|y���r���3?�,��i���,Bnƛ;�@ш�-�aP�w=����U|�s˦�NN�C�r6S��dY}2��j٫����E�$��[T��Y�� O�����^�� ����?�͊���i��;z��ݹ^��^S.�Г�������O��Szi��O�ҁ��),��K��I��"uU�\gw���@��û%X��2��6�z>nʍV�p���pD�{��*Z�U@q��d�M��l
HW�Tk�T9�o��1���BGf���s��&-#]B�O=g3���Riǟ���'R�Rc<H}�)eʀXC�������l����*��lG�\���Ck��'Y����u^��XNR�H~ﭢ��4����f�t笼�&S���T��Z��N�m�j�D�4���r�W�� ����9��]I!/�c�W�{��5��8)f/��-z������W���թ����H�ߚ�I_�$���0~�e���Ln���0|��������u�-�D�C�e1�u[�P6c/Σ��]�b;��pN��7x<�@����Ɠ�na�`�?���I-S4Z*��
��;>ُy�:����I�8��q���+��W"z��R�9�E9L�.ڂ���]��a����Y�dU���m�I|&���V���F>�1 z���|q@�@��d������+ݣ�f>z�Kv�!8!_О�k����yY0�Cn����'��B�J)ٟ7MH����_C��f��4$�|��3����w@�ƀة���}Y���DU$�+��Qˁ��p����>q!��#}rf���zb��C�	*��qݑD�C/\k>vX2R��	_���s�4��əM�<��h��<)J�&q�"�����g�V|�A�Տ��O]�2A�!e�~5��Q�!I*h����(ݷ���~	K���MS���0�D�7����Q&UC�&�o��3e�j��A��کRHJs��WJ-Rw`0�eM�ZV:�V�lF����:?�џH��60��v�q1_�cs.���XǇU2ӳ�%q�ft|�L��]�[�Zs6R]0��I���(���Cx�W%����A�h�6oh��"�W��gg�{y�q��P{c]
�ʞ���i���2£���Y����N�
�tjA�y��lׅ���T{�i��d�d"EP'"j��_7Q�t>�ކq�Ú6�WZ<e\0��U)k�$u��Q[ȱ��E�g��C~���+P1��ˍ-��|�zخ?M8����_����?]�����,��/S`�BMIw����aٿ=}��-@��"�pf��b� x��'oa��G�V�P��MUp��X�)���x˒p��/ӯ-�o�������L�ʵ>�1��yB�] �8A�z�̇'d��(�����'4pbMBkX�0���>�#�h�w$uZ�3Hvf9$����+��F+��eG�v��.ߪn~h|���c�4�O�;���-+2ؐԬ����`�=�A�a'�F�k�	<!�DH���·��$�����0�+��5�B��R��|��^7�C�6'y�������S_!͒�wZZ_	��G�^ 9��G.�A�pڌ�BB xO��Lv�H�gTR�'LXb���F��85w�	�0�,T7Ϧ���JH���=�;��8�_�v�����j��E5��+ʐф�ė��cq���UwC1� ,l����V�4���أ�9B�ʵ54�U�i������5L��d'����/�F�W����[�.\�Ayi͓��7
G\u�Rɖ��}����4cY��%ٗb��,~PH�H��@�_����eo$�L7!�5V�(�	x.4D�Z^Y����Ŕ�!��ÄPN8.yGj�n �"�T'���i��Άc����1Osb�z���g�1�kA�$�#�O-q�L�'
\z�U.��w�ݒ�48���Т��M:K/C�r�,8,Z��K���;�mWX���4��av����0�KCv��9^T�S�r��<dr���F�P#�FG�_��kҁ��ߧ�qIȦ��P�W�o���w�~�y�6	�R?�����`yx?4��m%;R������������÷��l%�@F2�\�Ft����9Sq2�}fD�.�Qg��(�¦��/�b8I�vޕ+�81�eے��<5�ӾJ`����-�[A�	{��/�j���_��m,�5'Z&)b΄��.�<%b�V9,�w`&*��v�N��@F���od8M����
���E����=��|�cĔb�#S�G��r�_�+pwJ8p��,%����;�.����]u�Ee�-k�{��6_�n�����E=��N</�����z�h�n*~�x�
�9��;��a8U���N�z�d�;��]+a'��l��۸�'�
�#3lڀ"Ct�*�n
�tO������q�2���+����<���-{��[ ڭ[7>����y��%^��Q��&; ����l���s�����z5�)+t����*9��[�NXs���|�|��<�
ט��-���c��	S��
{r$��ɾ���Pt���>��(�3���
B�%w/��mA��~2C�<�N�ͩR d����_;��y��/��`�,"X7f�gꥴ������.���O���k>�h�Y�٥i(��x��� ����2��,�P8���$�'6u=`���@�zTZ��y���4�x��K�;�����3�[�����q��l����J��;���qJ&�A0g���V.I���|Wׅ,�c�d�܌�]w���pG�y�a�1\Wr�P��_�(����u:���<�~�ya(=ŴE���uoٖ8��� f�雓һǏ��ܥ�謣�j�U��#Z���]+�I7G�I��>����sTS��<"�Sz�y��4i�D��[?ӈ���p�#�Lod6��?��+��k�t�`�gSKޱ�|nT�hӒp��;�`Д?qSD�~�	�S��er��^7cѬb--B�����A��}�I~Ig2{2\�ex#0_l��� ��P�<���0޸iMHD��L���9ٱ��s��u�������Fʮ*5da�_�g��d�ag]qLS :>�6�cA#>�X���[�f/0�H95�ih�n�uȿ8"ղC�M��8��2\�^Z��>�Mk3�X�W�lCz��q�I��AU��O��y{`�g�����6��@񙍳����?�'2�o�P�ʨ#�qf��N,� �d.�������)CWv`����k�θ��W%^1�H�F��G�7VףϙKV D��e�(�����$��}�����9CZ0���"�f���q�#��{`��}|��u��0��6����T�i����^�x���Pb�l�7+X_<�zIa��M��3�r8���J�:s�bG�O���Iy1��
Sݝ⼫ȶ/x�b�+��oaa�g %�*��zU��Q��Р4�~�}k�V{�&0��{��W(1���;[�*�2������$� �t����i��N�۩��Bm�s�����@��#�[��j��`&aQæ�:�yE��{�(��r� B��fV{���Is%�Z�b U���k�����R[����ʧ�����}A��SJ+���
�E�P���^\p:y2���l�j���T��f�P�B$������n�E�� �ߘh䒂�[�6m�({9���X���n���ʭK:�A�����MU���{5����� �����gK���2K�O$+~7z�J>���g7�E�x\x�]I��8�t������_�uA�`Q�.gp�Q�ˆ59�7�PD=ؿ��·	PIs���W�p�bm���(����k	n6�Pq����"
g�dqg�b-$�k�]��y��@;�y�mx��Uʒ��Fv�>� %k���uʟ;�D�6�:�ɖp���ɭ��9�S쀥���ojcV��n�)=���0nF�D`�vbMͧZC��{����n��/�s��:��GC�����M�aHt�p����L���������gu�G� �h���Ķ֪90Y�!�h O���l_�k�5_l�O�Ӗė]��5x�Y�hC5�Q�e�`�b5�֔/���3��I������R'�lK��k�2&�2���0�'��)��!d5�<-�R��>�n��
'�)ļ��3x~A�b:�)�ʋ��a����DƸ���#ϕf* ��=v���@e���յ�&R���i�.99?/Ǆpnn��T��+��T���������7�5n[�$!�c$NÕ�_&է�om��5�N/�H���z3Ă�d�M�d���ΘZ6~.w�di��\�ۍ�KŝԷ���N!�*��=H��GU�3?�7���įt��X~�[�}Hf �w���w�\HDYM.ɬ�;�_�S~(R�y����,�(O�����(������Q
R�����Ii��gLec�:$1T_�t�`�����F@,3�Δ#}���fe�!�G�����қ��S��
�2�^)..�'{&��C�7R�QG8��A�"\M������{��bܴ,{,�~��a���c~c2Ã�S�ɺ�g��0�>07�]g-/��2�&��������:���"���'���.H�s+�& ����=�;-�8Q-�؃�������J���E���)Q�^�;�G��Z��2�'u���O��D����6Z5RxI*мD���~���,j��s� UUbh�)Z5*� at6@J�s}i�m�g�\��>O�! rp}��;x(c%�^B�� �;|��,?A3��	��sm��u��>}e��6&��Fk��S��5}�r�q����Z�� <Ǉ�gq[�`�RObp�7�鴝����1�x�0��x ���h�F����RX��I�7��������,����T/;,��Z�o����,/0hU<~�l���S�x���n��̚)����S;3.f�E'���?wn1u��s������"^���NF�U���<U�9�t �)��ޮ��K���ǳUs�~aD�kJ[ڠ'�DUL��,̢m_��0�Jw ��!����������▅���H/�䪚o���d_l-c����T�m㥽�M[����?J�.�`?�h����MTKUTC���ZO�%�|N��rJ�2>��{��S�q�9�yLz7�<Ŕ�ԫ�r̐��������r�y�o,y"����������a���tZRIa �%��xʈ�f_�OɲH��&����Cf*{$���t�r���+� W��y��!�\��0���2=j�ئ�_����g�w�hC�|�p�r/&<i���M���5I淒9��y��7�)\f5�7i�@+\n.�J���)��q)	<�!FG���ӫ��'t����f6�>���t��7K%/��m]}���}����z�2�ٺ��:֥%�1��~��)�{����P�4�8 �5M܌{لzǜ��|K�A��e��.L
(���A,f��8�n9(�*�0�G�����hmPv�z�Z}�H��T
u�o�������gqO��a���a�_L�����İ���}`�Ӄ�b{Q��TR��O�7[G`�+bQP� ���7���v�L�To��ؑ��>�ޅ��+�Ή���ht<ի�u$ �K���Dc'c��I#��J��v%e,Ҝ�j*ef���e��%M(�d7y��<��N����V[�x�tҼ��Q����r�@S� �+�єw�Ч35%��y� 4�5��l3���V������LR|+¨�k�(�N}!��~��UW�w��X����]ݚ��x��v"#ǭ�HLi�J	�Id� 8t5�%��b�/�J���B#����#��7�n ��C>
ِ���LNVߒ:Uy>)M���jVwol��t'�쨾�?����Vl���(:�q5��Uyh�
ڑ�*}���3�R�[aQ߉��Ѯ������Μ�ʄL��ɕ��"��!�d=�S�6m�]cax��N)]��[�eG�ľ� "u%��Vޅ�C<�TWq��߷�pf�q��*��������͕�����/P}���C�b��[��:VY1Z�F�w2S�q/K��-�����P�� �f�g�s�Y)h�Ӳ�֬��7�Y��Τ��Q�.��ݷt���0���S�HA�U�ynE�L����A����o�����|3�&6	P\�
��4*�v��_�c�Ky�gr�e��7ѳ�I�.��V���u��v��Dt�ب��s�ؤơſf�!��Z�LTE�����n�/��e�3Y�I�f���w��O��R^�3�-�4���}Þ�C�WŔ����H�\��;�0�7Z$gpэ���`���
�b�~�̎�����aeI�;�&H�*�b���?wf�ĳ�4-c���@tb��ۇ2��*���ў�DW�9�H��:�Z���`��4
k��*a��b��o�8��Pu���{�o9c���27ʷ_B���6øQ&��k�s�?ٿbZY�̷Z�S���9��M��\��6��6gK��Ȟ\��)�G�����H��ڻ�[<�IS[kp�thS��ݡ�̥[��!��:�D��J*��֢�X>as����6�dZXm����;��	HceNÙ���Z�k�J����JV��C�\��	k�^S�8 �B�.ơӛ�	8R����4�B�Ip��i2�:mH���5=��j�ا*<�5x���_lex�y�!段��o�Q��>����� ~�ɻ��1�ݼ�=;��B].�3�Vq�yJ���,�;��-�ʹW�e�4d}�f��d"�a������5ƚp��4���~R�����&[~�34U�s�H���W�jh���b8٣���ۍ'�Pͪ$�'�K���#��#�
V*'C������fH"=���X�I�?-z�nJKg��Y>Ȥ>=�{6v���7pjs�f7Qt���&� ��LF��b��K3��!ln�pˊ�ਉ�-7۸彏F���C�=�����W�K2�u��N��h��VY�J�`����B億0M�4��&]ξ
;��$6q*�z�ʖZ��H+&�����σ��iox{�y?�mݣ�Ă�ڬ6���\o��I� y�	�Eţh�Z���BI����У��?�e�� T�my�C) j�i�C%d�m�[H� ^�4v���1�����,[Ŕ;E%�tc�o���h�^�����6�p�,]O�P�	��2�=%a�c�E�/OX������ސ���A���{q.�VA7��?��f�Fe�+̥F=��>����H�0)Į�`���l�o>�D�C54.�0$Q��߮���VM���B�=hw<�N���'����$7L2�
mGH5W�w���&"B�E�	{k_�"~��k�)̮�'/����W{~�[~8 �.��Wd>���S�H1�4�])4>�1���	; �����
Sa^��������qZt��S�K�Gq��f2�@7���td����sݢs���)�+%��$$Rl��J��#r\(��5�Kjj՛��XƤ�T^�a��s`Co�N��/[K-��e����8�\�$1V���1OU�g�b~���6���?�^�r/+/,�[]���ڼt��\����V���>��'G��`��w@S~uۭ���MM�lP�7�,��C	�~+b뼔�ؘ4����N��r��^@��Jy���%�"�f��^X�����i`��ŊKG���_7s�@E��:r���WAWI��8��M�b�xe�.^��2�j�qi��j��Zx��U�2y��0�
�m�^���5N�X�V@]��=�5��0��z��!�^q��7 ����餶�lw*���eHgr�������@�ti��U���#�-t�PZ���W��kI'�n�M_�?T����cڨ�-\�q���Cg��(Y�r��F!Z���� 0�}��=��ˁ�ڞÊ�W/�ߩY��'K��R�d�<J7��q	��f{a�`�N��րP�Oӝ�` �.T���E�M�T�S��<!=ӡ�F��M`�J��ƴ��4}Ĥ�ztQr���mԇ����?E')�ޡZB�*�\*r�� �5eJ�X�I���c�t�휷�O�U!�+�\S��_�Ee�d'V���ߘ� �(|[@g�$kS5�5�E4�����YF��B�v��{��]Nq�ި�9��L�#�kȚ0N��fE��E�᪂��EKL��d^�>�o��"��u���& \r��?�&5��&�x��,3��y��E��=r0[)��#�қA21)�D�k�?�&{=��fa���V����H@��n-����-70��S�+�R�z��pS��s���"1*���1ύ���VH�|�پ�?Yˮ�6_]�S�E�ͥ��m�c���
��{b�t9e��E��ư��:^c����Ю���㾋�$-��HA�����M�¹˘�<�\����u���d&F��iGsR��Ɇ5��F$GZG��2�^ְRr'f{,��6w��t ^$���<$wo6� 6�,�sQ&�Q9o��L�{Et�/����U�C�����!��|G5�3�Up�D�e�V��F<�\qծ��Hw������=e	!���rƮ�Don/�:�	�nٸ@�4�5��^R��Jٿ��B���·�Kex|~/a�Z(��ꊗ�_7<*�@�n0��g�7t�vS³\r�.��]�.����E�s��1B+�_J'�-���s�ʆ=��d����W�m_�5Y�L�E�\���j��t�)*�������Р����,#s}���������r�0���l.��
s�;�W�C���g]Srt�RRU�]�i�ǱIO�2$�j$�Iia�$�Z�3�q�	�5U"�za���:\��r���b��.��E�0΀�{A���+��/n*�һ
[C���u���@ʍ��g����w�˓����Q�Tp��C�騶�[��J��5��=����ėd���j��6�����P�r��� �iG\\N5�C�8^�	$����0�p�M[<�\����S�OCb�H���2�@�,?`s��E-i&ǿ�x���H����T�P����f�7-L&CF��U��W6|�/;�|���(�~{H<��8�:�5+.3��Y1^�s�Ɂ�o(4�1t-������^a����K��r����ו�����qض��?c���c��?8�#��e>�M :�o7�zK�(�7_�Њ���=˸b]�l�T?�P����w�{�HP�B�SKg�=TB�B��5�O��VH
��:�I���({�f��ó�:G��A����g8�hi�կ�0�"��
oX�d�l;��<[�i�=������D!�}]%��d��S����rbC�����y��Ȧg@n�k%�C�׽t��vK �1Uώ��ቍ�'��D�ԝ�
���b����9���Q�H�͏���Zi+��hA��_��t���3��F�e�-[k&����>�S.���XP����'�������eK��,�D��1V�Jݶ�c����jws5�P"��į�G�O���,&��l�.��e�-	�h��������-������S���$�􃵼2'����f��M�۫�)7�7����☎�*s�����3�pYζ�1�#"֠��Kޗ ˍ���K+���<��m��2���}�	���z�7F�WQ�2�~TQCH
�k�ƧV�Jyݫ�Չ��U��;��`%yg����i�K��`
�`8���cs �`I=���`��I{V�h|T��UIV������p2���V�a��'��aR��W�6xt/7��A���o��#��&;!ͦ�F��a��5����
�S�f(�b�E�I���/"ہB뙋��d&B#�I͡��PaJ���!�2�"�J�\�a�2�]��ӊA4&L�ZQ.��%�8�H��}:�#��?��^��W�(z=l�7:I��9��.����J��-lW�4���=�(�����D�-�z=w\g�M�,�N��P�_���ڔ���*&S��4��8��\4>0U�7Pꈯ|>MI��N�����Ê,9�y��5˾�x,�δ�`����=d�� �̓-z%+�1�4�4�����+K���|r���օ�:���0����T���Z�FQƶ��s�rQ4����4=Ti�t�!]F�E����_�f����=�Q��t'�Զ��bj��.ҙ�ߴ^W�0T�"��s�[���I��Ԓ�@�-��	��'*����}0>���ճ�*=��&"@�]0U����ŕ<��4 x��+��Z��<�&Y�#��K��!&U�?iPcrU��Nws��+�9�Hk��`[o#s������ʫ�r0̧S�y�"��:���",,[�5@�����b��=yf�(d�nQ�سߎ4��Y-D�6�5��:Qز�igO����="��a�w�5�N�.���ut�R�YW"�߳;�(6�S�������Fg��6g�c���y��NV��Tr�!�5k�ZWj���NK-Q~at��JcWk҇i�wn��|3���&z�8:�˿�O��a���7F�L�T+��G]�)�/,���j�d�!���lC�h��?������ڰ��#*��S���A������q:=8�(
(ϋ�yI�ț'��%�>BA�2�!h?�������D,�Y�_Ĺ�����5�E��Wr/'N���5hӒ��w{�j����^ S��w� !�F�c��MALm�G$7sx
L.�C�vs�|ri��(��0ф1�����6y^s]�)s�U,�41�^G��k�ޣu�N6��B�*T̥�=N��R�O������մ�GZ�>i>��=3ɍ���En��U���(7v�(S���ZM���@2�%]��Z#���
��T W�ci⍔�Zּlx��Z/�J��f�!9���'%�)yfw/Cx�tJ�5c!�,���*��s$x���B:u�+���J���\.e�P}� ����+�A��� �%[ֱph�U�	viʝ���Hn<z�M��9w�#��W1ʹ{I�H����G�R���3���0��~:a������r�x��it�>��\p���t0y�F�G5�:�D��>�I��B���$�k4�C���U����P$��3X���:}�~62~��_�X��M�V�b�v֟? <�H�j?�ȷ7n��c���&!�<s�e���i<�(+��y<��N�����1��4{C�D��p���Ggz�l���D���nZ��U����]꣰-��}ˏL�U|�+CIP�>X]5 �FI��vn~|�e�.Q�|M\�3�DF�AplZR7�o�9J��\I���"��n����I�Y�R��(33W+>A:q��$��W��4��i���H��vމ�3�3�O�ZQ�0'Co�D���>H�[l����̒ѾI�ږ��.��+΂�]��~����63űa�
�A���_��5�����O)5�j�鴗�����{CK�MN���1���d@e���k�xQxz�ŏ�h{������W:Ҵ(���vK�`A�J^k��Y 2�Ek@;�a���h:�-}=��v(:�`}�� ���L�"L�4����;�+������Q2^��&y�R�����z���l��(�uHH{�D{
��6�N��ui���Jk�D �ڄ�[��e�̀��O�oh�L�{���m�S�����]$ؤ�/�K=L���DAu��7����	���qe���?�Es\�ugV�3eL" ��k�Q�E�>)���ВL|�v����|���hd�((2zk�g�Te��WNt�`jgJ�[����u����nV.2��D��efC�Y��U�࿔�ѥAU?D�#�E��ʯ�n4�6rJ�N���Ks�?�j;�<�{g��РŰue�k�).��������6�/^K �Ⱦ`�^M��P��```�3J�w�>�w/�4���΂%| �����m��w⾠|�.��v"��s��ۘ#�*�D�~*�:AG[�d�1� �{g\���~��L|Ķ>�d�+ELdU�?A�zTh�ݗD9@g�(4HK%#�}.�~��nB\���gQ�T$x�p�]�)�o��w�I��O���,����rO�Z۽�� �g[��v�}�^pk��;�1:���p�6�z)@�F�����?#�'ʦ���şHz!��1%��CG9Iۧbՠ��aR�I�'O^��Myl��*�M���3�-���9��*3N]|�a��^��e!�����Y=�!��w�]�h��?f_���f�vRV��,��T�6H4W��q��xJ��Rx���-(�K���im�%%�%Z_���S.�Qϭtn}�2�2V��:(�ԁ&��P6C�����q2���m\L��iӴ��h	���4�!� ��E� vNb�T�����:Cd�Ǘ��N��2��\CSd	-�I�5��4��s=�.OvM��C�W��u�:��Ӿ8p��J؊W�t�-"�{|{�]��t�}%�7Srΰ&|��3'�H��k>��t�� ]���@�RIV�h�)�Ze%��L��z��&�:nb���zRR�_�t����x�-m�#פ�<��L ��q��K�ԉi��kØ�p�[��s�>��-�>t�9)'QJ@(��N��VF��xKK��I���I���	�d�+�F�tr��*��~�=W�'�W�nLo�ϻ��Ek:�^��$���`6h�G��tlF�����਒�:'��p5��%�}�a��o���Z���D�D��1	��V������߰��jfmM+�[��v���|��r�ӗ���
���Q�zrܴU�X�� L7�+M�����:��M�Yi�u4�,q~L��%��$�xe:��zlCZ�N�g�LJ�&F�6�#<�Z����fTq��6]�U���V"��mO\�e�&�֑Y!Ѩ�M�Z%��	Aa����Ģ������*Uܫ�4�h�s1�5�J9��& ,pSK��"4�TQ�][�4�b��h��j����;��V3��*���(+����<�b�=R�s���o�8�&�K9$��W��%�cA�ڄ^
d��X���HTL����>U�¤ ��7�wv�^��f�$�۳A4�$\��
=��K�,n.d����b���h��� IJ���x�7v��9���Q2�X3H5���&��mi(N����w�=�r�g�(�;����K�h�ȴ��9����)��+�q����\]0�o#>��#W�/.؛��'��Kf �	�G�U�}Z�0�x��soSxZ�p�(��]��+��$�al�)�f���F}�m�f~df�*hCZ��ѣ)��^��l��?�#�P�������N�r��|c����IK�������9
�B�#���Z"խe���A�ji.��5�nۓ���)����Ҁg�~�Id�#����4��|6���BT�:�^�}�7`l��t��an���JVv�K� �{�6���?�hl�wk��l�Ǜ�tQ@��e�<j�|��9�;H+1�Tʴg]���歊���:����&�ܳ9�l ���rlQ�T�ށ�p?��ؚ�zX~G�t�X�M�Z(��Onx�"��`����-'�fz\7P��ae�p �( '(�@�!InS��r(�hC:Y҅_l�����-PB{�pz��k�AL���N`٪l`{ >8$+�B�ڀ�9��Yz^��ž�|��l�o�yp��; ~R[��=H̪�Q��U=4�	��k���[�8{����ƄW�R?(�`|�Bs�w��bT�̭�A�۠h屿�FAf��{����~&�a�G�-��ZLx ���e������`�aG; �1�
xnl�Y��^�'�Y��a��p�1��/eZ�	�l��U	���+U-Fm?<
'}�����L	Jؾ�0�{Ooz�0��=CK��X�G�륙,v��Vt@M�`�ʢ!�"�p��8�9��|��xh�DuK��l��Q�p>�̚���� ���8�K4�k�De�/j��q�7��n���� ��n~@�ѿ����t=`�$xs%�����V��Iu%��;�}=�ù��A��â��-�=�!#VG<�<��`C������s�
��rpFs1�m6%?�H �<]�H!�6�3Ĺ�X���m�����x����\kwM�AՌc����c]����!��˛\TH��꽢�[��*c����a�GfKq5�zCO�$g����S��Ҙ:|5��ǁ�v�����ZҌ�/lk�N�xMD�����f$�P���BO�B~Ջ��S��j�*s�S�����ӷ�S8��M��)a���}B� 4���[����'5&8u�7)��,�٣V�4h�\�o`�X���,������K8��X����F�^�rZ�S�p���I)����Z��� � � +�+��!-�~�QvE�惗!uXzN҂�i��<hQ����xz��]��yF�QT�x�$+���J>�s:���ցF����������e5���j��Cͱ�����[T�R�<�Ĩcq�;��e<������uBR��3���S�8��J�:���#�Y��*t�A��[!m	����Ԣ��x)����%���_������up�M���鴶�x'��Wj9�T��/��{�y�MM1�Ѹc��0�ͨ.z�r%N���V��-%c.b�!S9a����Ƞ"��}mM��8�U���{�R�BxM0�QJ��Z��S�ˠ,�q�@s#�?��.I�3�(N���T��1n�Ti8Ч�:>���\J���0Cti����'�\�qܿ�z��|-B���4�����U���`��,A��1�a��n�<��x;�p/�7OYhI��C�J�݂�Ԓn;^��A)yj�d8 Mb� �a�ӗ�GAd]�������?o��ʞ@v�*T�r���v�����̽N�"y�L����`CLy�m����(��HqD��shNCtR�ʇ�ꖂ=}�{3�s�O���s����{�j��]������{�QC��V3�1��~-�Lv�p:��l��Й���~`4����Av]���;Fnh��9`)��O�.`Ř~֧
�uQ�d�]�%���,@{OExg
86���|{M �ܾ��C��}�.{����;J��k�����h6Q@V.���`r�e�}� ���]W�q�]x"$M��P��B��K�ΜA�����Q�E�������r>Ψ�O�42��C';(fk���������.!:�e�]�Ok���`#�˝��21�TȰA�_U_�*��Ed��.��h�
8�)�ҍ5�ő��v{���R����ڽ�vX�6�mOS�~��"����L(�#�$n|V�K�,������<��V�m�47!�\��3�s��Gd�FF���ڟm�`�F:*�w�gl4O���{?,?1�Q���f��.�(w�7�5b�6����$Nw��bi� ����ҕǧ��j�����u�U��iߋ��78�g���N��.���d甛�����D�\BJ�x8�i��5=���N���+*gv�{�6��*3B���\��kAh�U�FS��3̟ǩ�'��x�1��8ԓ�2��e}�+��W��Q?N"�B��&�<��Hΐ����U�-��]ظX	�'��9��$公aJ�h�p{�aR��v!\B�QL�2cTXV�S������������<`���`X�XH,��q���Q���R�=�a*�(�L.	����@1i�y���owy������H�v�p��'WLf�����m>�yj������I�z�-N�J>,����rج՘<��Y�ӿM��?u����km�^h����.��n�I��z
�gm[�� x��t�:�A�8�+��6�Տ����@�W�t�d]��/���#܅��U��i�#K"�������T����j|b�TR ��,�O�L�PG�"ǃُ���"w��j>�8��	����=.P��:%O�٣���g�~m� SE��z�� ����ˁbNX�l���<K�T����.]�_�Ц;BX���+sv�f����3�{M���JH�&.�~=�o�	A������?z#[�-�	�j�/��/(�rvMDֿ�pއ����Y�3 A<�*�OZ��g��6��{[��M�v\��U�f�x�ٌ��y7��آ{Y"lQ�'z��Bq�l1y����y�}5O�hۃk��	�crf�혦C��K���?y�ĻU>y&L5:V#�V�� ���׫)^�b�Z~��tk\��ρ��V�'��� hX!�x�[��E,��/F8}PZ�)l,�����Bm$~��ON^JF}U�񼫷��9?$�N:�߳�9�:+C/l-�!�զf�$�u�>�/M��uQ~��)U�Vh�9+"|V��x���)1�]I��
j�Z�=$���=�l����7�R���l$VU_� ������;U[=Y��[���8O���� ��&^�|�1P?�v+�P+P��Q�:��z��N��i	:����q2B��gy�ߐgޏX�?�����]�Տ�sp�Y3��<v�	�u�5�]�+������Ԥ_����e��k\�P-p|� ���J��BEQ9L��<%�P���D�m�����S"��(k�%1�2%�����Q�"h�q4�Z���ςau;��b%(c4�Z�1g���-(�'vXk�f����{�"vD�U��\��9/�rH�O;��E��0��A���d�f��8QmKO�d6�#Ɣa�c�3��A�Z�*��I����6�˹���H�y�ԥ��Qs^O�n�ZL5��-"l�o7��B��w����%�K3CL�l�̢���4l�;	bi���}�6ܰD�w��(�)��ÀW�-lv�#�}a,��H�W���+����3A�$a�&"�MV�u��~��p��(2������}�9���^N�`�Kb��o=��-��]�נ�ͿX���w*�;���H��Q޺�s��.�8X�����	��Ry)m�<k�0���"�a^� �B1DӡRMD740��� �c�Ԅ[���O�ӷ�߉_���܉��8��PvS�j���8J{'�I���`�6����j�4y����� ��q���[}�{	qR%M��Q���!I�uL�^�@���Wms��b��:�&M�.�qF����ں��eDc�Fj�Y�����=��ե���s��H!�I}�����p��/��$�����s��1���]u��X�+Z�(I��e���J�~fBlW��F궎�\蔵�l	�6<�a2�Mo�+�Lc�2aNI��afs�Kjқ�X[�$�����e����d+l
� r�k�l8K��@��NU6��Y�	xX:�{\��0��$��^��E�4=�H��J��}�"1zYɩS�� i���`�gVp^�H�b_AYK5�_X҃;�����DͪM&�as�L��4l��k��5콣2� R�<�%�.�>�`,����8�
�tX��6�ʎF�w�-�(ГI�M������*8�	�#!��z̶�h�c?΢|J ���)��j�L��,�'�ʬ�����5����b���d.cb�w�)*�N	�����T:'n0K��B�|6�!b`��|����}��)\���e����۔IH&bs/g�4ٴh\v[�d6�!e�������������~���t��.q���`f�)\���F���1gn6�={�h��%J�&�ѻ14����Uf�p�3ti�T���rEj(��6ӕ[2���ڧ��C�����H�U-2��Y���d٥z�q��{�.��+f������B&��M4��p�g�cßw��D�'���pq��[�O�1�pN�s/�KZ�lz����,�W��~}���[��E�*\�C�cϴ� Y���4쟳o2һ(�D*��������z���tjθr3T?�خw�z��������r"���ȳ%�Zb�3Ϸ7�3k_ddw{�1�� �"��Ӹɴ����"I��F�b�����oK������	D=�ȯ��t�����2	��c>�A�pvג����F���ھ=M������YN�r����U9��C����	��<�#N
㿼�כ5�x����L�֊o�E*�R�Z�tW��Bi���+�$�fX؎2��`��	�9�=-�*�֣�1�z+ގ2���?�2�!���������[�#��k܀r9��^������>��?v��XQ�i���FY�Q\.�ff�h��)X7J>��VR�/pZ�Ƶ���l����o�C1�b˚6�qs\m�J��W���p]�0u��j;���fx��jm�� ������ԨS��i�Ro���cD�?W6V�2x��:�O`Z�ܐ/��2���IOW�x�a�\�I@�3P�zQ����o$�j[�b$,�M(�-Pt��P��%pA����n��b�8ۜ~���<!�Ɗ���!V $�����D͍i��*���(�4~qrJ�M�R��>i��C�,e�ЍVG����X��!�>��kT@�_�=+D�n,Aر��!%�F&%���k-��O9��<oW��e�Rqd�{۩}rb�X�N�H�0����S��Ȣ`���ߔ�$��us�/����dQZG����9�
{uĮ������*�v%��{t,;�m��T��W��^D�S���u:�P����7�}�r�=���Oh�n������c�,s"|���|�ZbT���g�k^���D�>��u������El;�U8��TG<;gl��F�ᡈO�HiЇX��իr�H�K c�V2�X�Xqt��*[���!����]2�f���e�a5i�	
��f��VΗ�䜯Q}g�[RrG���'�:�Q�2%-¶Pm��Ug4H�������uJ=�*s�$�V���>�WI[��ɀ�0k���n&���J�z��/���.b<�K��-,)��O|CGY�m߅c���V���%�H��Q��X��ך�/9E�׬�9~�F����vPU�+	��W�C@_$�:-�/�G�:���6�E�+�E�\n!�
�y|�-)SN��� ݓ����}?�\��(p�r>Sq- �>7`�L�|X@tހ���?��F�iS׷���s���38�^��^&���u������;w��ep:�3e�t��^�A���[�tr��'�@еI���Wv1��~BSh@�[�Zϥ��})"zFz���ʱ�M�
p:�^G�5E��#�$���I�A���P���,��7�?C�#����\�=ϯ�K��!h�Õ۝�=�x{'��:"�/��T�c�Ɣ쇻��t����ޭ�d��ا��m���F%0��be�����$e����^��O�r��=>R���]Iz�]������1���s�͒�x.
͂/�{We�W?�����}��c@�����<�N��	��o�����(��u/%ۛ�h�a(KVU��a*Y���x� ����[�����+�i<&��S}�
P�X���	wqi�w��0��!�N�39} �[a
��y-�ٌ^p�.�c�Y�EY蠁c�nP9�4�k�����y'm����Il�!��`�g���/����n�����%in�DPT��wem�p���P����|b'�j��ț���>��f�TÁ��.:���`���)2QU��?�{�D*bS������L�b%	J��� �E��V<[�@.��o�(���M�՞��Mҩ��r�6�qO8�����EN��&���>/�%+�n��b��ET�J��`q�5=�R������V��x�ޥ�uo�Bn%�>MI��!�Ɇ�'d�8i\�i��"�6��i�*`�z��/�#��"�=���=�'��ۓ�x[,MRF,�	4w���x�3��%���e��_7��S�Q�4�Լ÷�{�KuH^��̲3��X��io6��w����b\0�B#��yZ�0]Rm"�r��y��юሤ63\�w:Y;$��'<��*|�{�-B)�!��I��?�%kˠ��j��p&�f��U��"C����i����Mh�'�l4��f����{�Ĺ�ĉ�kDlQ�|fB���O�ԥG�ȃ�V�1�p�I�j*�b��
�@����ԙD������m���c-�6.\[Z�NNƤTkeCre�4����ѯ@�jm��{*Y7�G��i�TE̱!J�U,�)����H�M(M�/�I/�u����d(�
���\pU�s���Bٟ7FM��{C����6s$s��(�j
n�&\Ef��]x�[-~��ZHFU�K׫���X�{�����7�?z����V�w�.a��Q�
l̻��ڔG���Tz������-I�0�����4���r��,��M^i@m������"���2Ϯ���˹p6�p���K&%���g�����y��y�?
�_)� G)��`��zs�Ϊ0��}�_�2���ʓ�������W�d�suX�������'��3�u󑯐�����F�����@"d�!l����nm�,t�o�>���U��Er�{���A��
 E��Vy�H���xmw`а�	}�}�e�2F~͒�e$C$vd�օ�#�� �sNd4���r�/ ���ڟ�ǧ�co̜pL�T��Q�:�F�c2���ydX��1+�>�W���7o��T�׍s�����#1�;5r�L�js�f;ܳd��Szs/K�%Q]̲�����:�6�e縘Y�l�2ū�͵<I5 eO�r���uX����B��.h��{!yA�Hٻy�����fQLy��Jk�6)�m�=�� �Ol�8ɄP`kG�#<���\��������԰�p����~��+j�y�Z��d�r���\7�6jF�>��9������2�x'�<_��#�7#ML��5����9�h{]������ÿ�$$e�QטE�ּ�:��Պ��"�DE��c7�g^�nPf���~e�va�KV�z��j�f��A��)���4� m��ך]�>�W�͇�[������4�>o�����O*m�ke�[QR%��`/�M�Sݤ]+�Nф��J�\Ȟ{fh�g!��2�ކ�B�e�/d)���Aܔ�,�YrO�����#r�Hf����]Wr�̵m�N�Zu�J>�]�]����c���n&�g�x���2mf��gr03WX�6��F���X�#���]�5�ϩ��b�@\���+�u��=^�|��g���E�٘��G[�7�|bB'W���%���2{���y/��ܕqRVB	A�m��� ������%�q[ș�t�X�W��J��M�R�ܳ93�=	>}�a`��B�[k�?0�d�hwqc��nn-Op��Z9n��=��3CZFpq�x���j��A�n��Z�^�n^k�^Y>�':@?�[ �TT�?l�y�IP��i㜅��CN	��۾tGe'd9\���g�T��Ƨ��-3�dÿy ը&��xO�s�Bi)XOT���e%^��Š�̖$d'7"+P�����d�I�b�$���B��-��|�0��Vo9�?)�Kb|ȻK���]�D,"ՠ+�{��{��I�a�K6����l?M!q���?�(~�R��#D���T-�n�s���ٞ�#�4~Ӓg����)O���$%fBԊ-~R�E��u�Ԉ����Ȍs��n�Keh�f�l���9�\���D�S�k�R��;_+��S�c�з��).c���;�X˘�c�G��Ӥ�g��U��� 6�����6��8i�"�V�~&q�� �(�,@3����%�#}s��%"y�S�N�~-r��!
�B\�C�o(N@=;��i@�z�Hm#0�"�,M�n���fE�͟����n�2�Ô���D믲�� qF�F�ѭ�"p�9i���|c�'j������^^C�����3@c������A��mq؉}�j��$��=���>�˳���J��T/�bJ�H���IS?[p�VƭK����4������8�!e/jo��6~ugc��M��e-�Vxʻ�Br(�M��O6hV؋?
��UǗz��?;��9�5�����RH���C!�uXb�M#}6��L|������h�����GT����K]@�(M?��z�.�H���.I(���n珼̫^U�yc��RU�ܜ��¡�i�;��Gd�5_���G�`�����<m(^�?Pa�P��N�����>�-�5xP�a������Q2-�9��}fk8��-汨�Pأ�D����GB5��E���dB
��8x��_/MmMZD<��kO��������`䪖�+�F��:=�Ez;0��tb�2�	
��Fs#H�UO��`�3:U'1���xUA0~̞w��>� ���]�3"�gp�]k�8���>�9n���aBx��Φ�=G}/�?j͢"��JPT�m�'�Q�#�Tz���6��p9ջ&d;�aThQ*�dr"�U�8�Lg)?���Y=.�:~0U)�:�>f��KĪ�WU�Q�~O��=˹�R��D-�ɥ����K�w�(�S�N���B~�ܾio8��0�9�S���U(���E'��7��^_v^/����p�V�kU����o�I��, ���Yo�a��Fp�鿾�YU����Ւ�c%,��;�}�%�$�*k|o�Q;B�M5/���AA�; S*���\4U�)���$�o3��k�2�St W[�C<@:k�y�n�$��{��YxV9h��ܖU�0�(�C��QӴ�]�=����bC]�������D��}(���}5e����g�����6�/-�@��,�J�E ��$E�킟Ѡ=E��"�w��$de����)bd�|$��]z�l�cT����Y�'��#V��B�'}�c�J�0�`C��������W��s�����;8$�͚���"v�|�{#��`�c�M(8�Xk�u�O��k1&xE硶�1�k;���78 �"���rF1�S,��=&u�va����6���wՎB�Y;�{=�^��q��*~�V�/g�$S��4 <'����;l�,B�O�7Q��Eb$�q�sX���֠*T���Q.vQ�����w�:���9M��Q&JW0_�Ex%䛙;u ��P=6�G��pvI�պ�6�3�όD�[ -�ZIZk��v �5:v%h>R�o�0�@��Y}_�wk������6�ԥ}����ۈ�${"�@N������>�����?�+�,�-�:����J�Λ8�D�ܒ��/K��7�+�-����8W5|�el�`q����T0Ǽfṋ#`�r��&�"�t�-:Y���2��I���,������0�-d��C0�(������NOl^���y7R
ܶjI&��G�M� '��XD�-*	���1b֭$����l}�.�Ք����w��Z��%1��ϔ�ȍa�q@Bߏg�]�\��a��՗�tOs ���"�G�y�ԽՉ�]{.�u��#�����"x|h�<������q���D���`+)�_�� r��F�UU�z��D��RQ;b�ԛ�]��D�*k��nS�̂���?:��s�'ԝSk���Sx�-=�.�G�	��DK�Ѡ)���O���ʆ�NT�Y�]a�e\6r�|�.�Ki��B�H�e�?ag����qֽ�0�W�ܦ��q+�,�lo(�5�P��]��@�%�"����K�G�d2u�0M��-�M��wN��=�vW	D�$!���{G���%Ёn�d����R�c�G��ȹ����:'[k6��ӧ���2��Y��WWQ�7�n{WiBj�n�`۩�^�0�Pa�Ҭv�G��E
�sM=��WKF���C;���C/�����=?u���~�@b��D��FN����ɖ�X�H� r՗�1_i��ȯ��e�Q�/QZ�z�3�Bg����ꖑ�Z�>����kH�q����1�ÛR��{����G�VA�c�@PLq�7Y�N8	�����w]L�/���l�̫$�\�X��E�p��)�#��ō#ڱG��$.Ʈ&�/	cn�Uw5(B{�~���+����q��UD�����
�T5Ж�n����u�~�D���pg�~���=�K���Q@寰s.�V����zKx���$}�K<�j��͌b������n�X5_��%��y3xOݖ�{4�h�=�����^�g��WoC~����.9����E�l��+��D9J5�Y6s���pȲB����
Ƅ��/����BK9<=��s�0'���7�v/ȶK����L7���5�>d���>q��R���:;�[�⊔+�[�D�����^I���x���1Y�i���D�S=Z����cٹ�	?"�D�#�R� �jh����y[��Dz#��֜Z�T;�C��"�:�IM�|����?��B�1����_Ȃl;M
�w��<\��=�M~�ee��Ps��<��A����i���r���3�[����U/��=��ɓν��2���=>����1�W_��$�0�q�C�&�����9S�%_��rS�%H���zb@���>hFL  � �ܒ"����}8ty+�p@o��K��p-��{�[�H�H��W��H5�x[�qO�w�Ft`	V>x-4.���/+��3k�PZ^y� �J�9���#៌���sdD��ޤA��W�3[�c���db�%xT�:��������.5��dS^
2)7<"��k��C��Q)Y��LA?a�}y�]"��3kB쥳�]7�p�en�x���\�]X��Pt|��Ԙ\k]��!������8ay`���]�j<:�ϞK�>? �|�����2'%+o	�(Y&-]��H�#km�s��$���8��D `n
-�O�}VXqU%�V	���w܍�5܍�A����B�2��xGH+�,�x���S�>JĶ�{պ�pA���U��}�3���^%ޏB����WwF[���d ���ZH3#�Y8�3��i����a�( �
ېB�@?;��<��*�(�n1�� l���0�um,:޽��+��Ǳ�Ǝ[�p����MEkj���L�T�:,̎�gl`+������I�&�����ffyx׈C����BA?��	���/X��c��$wg2T9'�r��}�iʹ�D~�k�U�����zG�W������-����M�����!��[�O\�83��c[�0Gg^i,�U�5A� MH|y��g^�v_�)͓q"(�H��K��(;h0�W�^��Ɩ&8u�u�6O6|�=r��{V����b�m��R���oN��T+%%���X�<��f�Ȗ"���@�-PL�~v��\�՘}�hS�SS�� 
͗T�J[]o^�^�p��.e/m>ڌ��}�� ���&��tx�>)��OU)�g�>
���'g�bƾѸ�N��L��D }J|��2��{�MH^ƻ��$m�v���|�YߊmЬױ�]�S��&�%{WML��vH�da�-U&vP����Vw�#���Ҙ�5�U�3�;{�nT�� ��}�����R�2�X�!�0��4��W��V`ЖL�dO�j�\��9w�U Y��{K��5`^[P{���u�*M��$��݊��ZD�^�/m4aqF&�M�i���Q� ��(L1A�PF�_�Z�������;�fU��X�<�2**Z%��$!a�!P�V�qRGȚspq%�|���!�oPP����z`�'L,=�>CpHb"d!c�?�*��Pr�sL�꼁%e�T F�S�y�3Gߑ
R̐A�vAd�pˇ!��B��~�w�s��C�AԉCש� �B�7���i�&��,���K��:��c�2�D(���@R>)2/�:eW��4���7��:����$�'#}�9�|��Q���X����^���(�a��*��� ��8o�PK5Z��|r�\����p(���?Z:U`��e��m�W�'�����;��r��QP�ؒ@�}q5s�r�16���uT�沿��0���mJSc�P^C:���|�駸;�Φ���ʘIy2;�PJ��9� e���(�م��i���B���Ĝ:���ɬU����Ԕ��^�_XO�+���K����4��[5�	=\�d������(��82=V���Y[�5�\������"H��I��Xh�bk��_I���ԛ�PI^�H�,�A�R��|!p�.�R�Domw������i��BII�
��4�O�.C!N�I�ֶ�핸H֑X*���[��+B�d��F�.�0�w?��{ǥ���v�Iڍ�P�<:��>h������J���,u��ǸC݅3��6m��w�-�׋f������h��z>2�4�c�*��:$� ��;�E-V�|���S��������E@v�xR>(qt�sX��?�i`ZyY�v�F8�G�q'WF�]�2��x_������VGhb��aV�;���MߡG]�U���-b��{J�,�P��d�4��%��+�ئ��}�����������̧�_���9�e�N`��K��l�>�)gx��L��|m���;��&6G�G�v8
�!���>يޗ�$ ���'��AGD�O�2���!l3+S(2����W���?���)}��%�#j��7B���[À�*���4��,UT�iy+ZZ���y�Y�,|pa���"וҮ9��G�XZ�|L���QK���#h��!�0�8�'�H���l��(1{�uy'��4
V�'?��������;|��<!�����!�Y"*t�'U�mdky��OhQ�#
���� ���^�`�*���3g2�5"�`�E��3�݂���QjA��g����,��	�&j]#�����7z���U��ؖRI�FK$�����-���H��A�pU���R�#)�we�� q.|���m�����e��癩t��K����*AY<(y/^�ޑ�&�� �@>�H�f��r���}�A����.�Q1���B8�N�����X��� /M#bE�����d�O�:^:��dxk=O�/c�1�K��"t%�ˆ~G+aF\!V�����oz2�N��c�	E&�)V����-�l澆��5�0!��z��]x�)���]4�ژA�~����I�쳟m�)=e)�`�kl�ʋP�P��Y�w?����f!h垓轾սe���h�J��{�^�	��rp,�m3�<�L�5�:zBz[źL����{ �����b�y�|\�����޾r`||�������ˀc�[�\P�Vs|x��@�9���a�,�"{�Y����+�D�%��g�����p�Z���	��1��`�ߚ��eP���#M�ɷ���q�uH��R� `��oP�;f�t<1���#����\RR8y�����m���O[��-2Y�]��N�txv�O��ڍ���I����i�D������kjm�Y���!W�e�}4Q����EI�d���u2�ok�b�!y��,�(����B�v\���`�e���)�������۞/�N�q�8��7"�
"_�p�b;����uȄ�W����[u0C��8�^R�T>��=[�'&z!B�A�O15Q�Yt�Kz�L�(���0I�D�e���J�� ���耮$��8�-s����R�N�:� �W}�0~���n`�B��O�=Q�E���u�-s���?Dl�����׏�9�j�0�N�ӠK5��IQҢ� �rٞ����p2[�ޞ��(i�(н��u�iy_l8���01#
�l!mj=[ ]�܍ۿ?)�*�'#������3aںy\D&���N��S�������=;��KzS	G���F\!v6�/����Z5� ���u@c}W���u3��׮E���.;�]8#����]NN}��B~j���K�vuA�����`�ر��-�����(���ׁu����Cxd��� �#c͙�������h�T��5�mlS�f �L�2u����
����c���{�Whl�B��$�ʱ���,��=��r�Ս�=��5G�4K��,J�������,9��-�p�'t�Unqq/��*��v]����g=�^���	��~R*6Oх|/] t�dN�&!��0c������R��+މ�C���w�Foޚ`gs����`b�=t�5	(��������R��!�Ћ��|Rm�*N�sNW;�SP�jQ݉��kowi���{HD���4e�h�JC����l�o=�%������xٚ�{���K �K�R�K0�JFcΒ\_b\�1�p)xk���@Y�`�~�4�6;r�w�&ԓ����a	�%�ᎂ+4�'pY>�j^�wM�E�����S-y9^l�����f�X�O4�j	�a�qW@�Ә����XP��y��	yG��M+����n�Q[�xڒǌ�˭�~`��o��d[[!}�p��!�@��0>BN|)��x���� �9�
03�ȏ3+��Y�S\C�Q:�V��R%��زkZ:*�) T���JC�E�=bU���t�N���4�������Rn(�&+�O�� ��3M�������pwp��jR�e|�֊xvAm�>�L`t�6[��EH�'݉���l������>\?�\4��-�؁���~!�_v�ӱD��Pi:���֕�%�Ys�Q�I�<������?)��z�x.����-��e���V����T9Wm�T��*�x�������yoJW��GI@�cL���a(�<����j_��_��F~��7r�Zħ�sWf���߬}x�q�r6�Pc+@�v�jc9���tƇ�lϷ���O�jk���s�b.���3#K�K���&���� 2D�s"` E�ll�w�S|�{X9G;����>pH��!zjQjGx��
wi%�e���:���zAu�SY����������͸���&`��ڇ�IWM]��[t?p�y�5p��+
y�,¦�����-�	���\����m#E���Ovj=)zK>>�Fj�R�%���O�X���|>0���o��8pz���7��To�%Ƹ���ԭ�i�V8�?��h������\���7)-t
�z�)�d,O]u;��y�h����Y+��K�O�A,�^߯��V+�w3G���SV9����b�kc�}f˗�U'�H@��^[��A��m�O:�G�� w�{�D�ei�H�Lɭ͙�u2�O�ޮzᅙ��)(��<`[&8�������C���pR���2��$���]���O�5x�?�}'΢XWgͶ-��k�����̉�������j*���=7�.��B�6�s؍��OA�FGt�N�[N����cf�Pt��5�d�x�9Q��񇣟P"��3��v�I@!MZ')k�x�i5=��f���UkiE�<%�(�-h0�g�f0������`M˥W��¡��64D�y�44e�b"���ΖYHH��ǯ�纍��}�'�8���Ɏ��Z��+�aw\I���:Ay,C%Z�.|�m�5G����᪊9�
�K�M<�]�����#����T)�*���DsX��?�}tp~�{aPbvZ}���*��O�ˈz@g�(�5Ayj�ț��ft�G�d�H�� TJ9��s��JH1@��bX�|q	�*����d$�� ���в��A�R@��:�盬r�l�eX��2XLfT�Cϸh��PQ��,I�6�s���鯥�`V���9*yɥ�D�q�;��^�Tg,�<��n&�z�V���[��l��l�O]&DH6!���(��m�>���CL��	G���R"�}o�)۱�Ê�������
��$��\��Mv}��/����7S��j��cQ�(��z�kK��|�B�%^����QUzO���v�`O)Z�~d�������P���u|�Ӟ�z2�k*lqh:��V�n�X��Mø2�Zp�dt"2�LP�-����F�p��h��.¹�w���s���r^�4�i$���Z�9����<�Vt節��N�q��ct�O��+�T��g8��"y>��_±�t�����szu�`�)�G[?m4�,�e���_Z�KT�t�-�iu�FH4یܕ���� ~�T��� p�D�������z�|�["EƩi��&���:�����e��,�856� <i-�5��i>�\�I5k B/s��p��}��n���D��
��[��+���@�,��х� ��t���ꤟQV��@�jNA��?;�+����4?C�eX�]�V)�0+ ����D[�t�]���Ѣ#������0��m�`>u�" ����^���d>r�{�[!���"p�oN����6Y85�AJ�E�$;è�s�.^��՝V�	��}�U�)�䀹��/��w� $��#�0�DU^��>��������żK=�4f��@rX�5�v�}�;H��Ņ^��O#쇠G���:N5P$_Y}��*Zζ�*�W�%��l�y�j>�Ң�����h��u��=S1(>z[r���n�s�r坫{���P?�z6G㼬� �����x�B@��zCx��g�hy�l�z#tKa��F��x%��z. ��R3�)%~�����f�`8)��(��g��F�\�v,3Y�Ѣ��?�;-�-�;�u�a�?�vG��T�$��LV���&]n��Tq떫1;(�8����."���T@w]TG� �9.
�>�����A2�A%[v��5�^6���Ԭ�-�~X����y�B�X[Q����4y��Wy�������=�7�+0=N%��`�+x�Nc]��y��4��q��ߊ ݗ�}Ab������︐�kN���Q��	�%z�L��)�|��kB��٧qӇ�B/�](n�L�Rňϧ
-�o���<9i���u]LD�n��eͣ&�/	�Q�N
^&�Q*;��ɒh_���r�\6���	�Ѯ�Sן���4Ғu��0��)�IΦ���T���Ɋ�m��R�4V �ic��|�y�\q�Ң<��Ѩ#!i~d�{Ʋ��~} U"�6Fa�/����l���ہ���c3t˾���a�J7;�>?��\:����m~5
����'���Ƙ��V�b��+/A����[�z�����k׏-B��=���j/'�"t#q�n�>�!��ɏ��C`7�KQ��e4��@ �&��'m�VG��w�Ϸ�S)ˮW�Ig�5LGl�'��=t�H)�P'�P?�^�-�S$��R�4=�`֊#x���o	�e�c���ξpZ��o��, @�j]��6s�_h���f����d7��uf	.�i��&��$��ߜ�Tb���Ob�$���w�Cќ/B���#3o	��e��D|�uc��$9sx>�'M��S),Q�����W>�<��Z[Ѻ�
�Z����l�ȩ�� ��8�!��*{� �`�ر�,0�j�6�2}� ���	�I]��fo��Uue������>���>H�*��ޜ�R��կ�kn�Y����J��<h/!~�aY�A�P�����б2�Q\����g�>2%}["�g5�n�����9vw5�z���)�삶K�{ ��X��h�^�;+V߿/��2O�a�!����٥'���Z駯�\�g�_T���/��P����M8���7X7V���|����Q�d�`W�ުȨ�z���4*pSwZNMv����H�ީ�n0���
�w�.c�A�����~'P�9sw��Ղ�Е߹6��Y��\����K���k{(�.����ѯ1\հzx慊<����'a��&�hy>uI��u&٠5!�� u�.���U��rƳ�n�WΥ���u{8Z������c���ڜ�-�5��� ���%)�9�������{�,n5��Ɩ1�b����X����5�� ��PYRW�;m��$|W�m@mMc1�z��F�_�J��.;~\��!��S".�7���^�6���C���}=��S�3H鋑'�Z�	�)�BT�i�e�s�7�M���zD47�N,�%�|�[[_���y���	�+�t�6/ާ�A&�w�~�/&]�n�������(M?w,>_J�Ӓ����q�6�� S|k|��_	�T�*tl�Z����E�]ħ����;�y���<h�k��c��%
���´Pv4ⰵ� �u�(���,9�C���� )�X�
9��b��6zD30j��^�7�|9�����WA6W��t����;=���](����[&��A�{T�U��?ɀ�N�V���C�� (���(��i��vT�g~&�B��s�rs�V�%��	.lW��(5Fϥ�kw��!�q�e�
�{|�E��G�t��9�"7Pt�ᤇ�ڱȵ���\��P�$�^�0�ï�>LϮC�#;F�#O��[��)���� ���������mq�,g?��mk�*f�Xo���qh�,���Ec��?
�!��q�1�,}����T?��2�p�O�k��x#>���a��2�A�1�b�y)b�|z���
�*@��}x%|t�͆��1�4C��c��u�A5��2� �qa0\i�r��@�$����~���!�f؆ɵ�;v��j��,5�ܽO|涀0,�}N�M��B�bQAm��B(MZ���.1�� @GҡQV5$NS�TA/�z��}Kt���U�>�r���ӆj+��Z'����GèUc�����.l7��;�P��d,ľ+آ�j��n9@�EK�䓴4�k�}�B�*(�<,������>jMQ�,)VLy���_B����:Ja��X���Y�:�5H�Y��Ƥ��T�fbp��3GE7>�꿖�Ub�dʉ�hX@j��3�8�=��΅"�|3��=P��{w�����
ް�9��H�!^��W��'/r�d� ���)��PDi���{1MQ����ĸb7]��?v���u���/_���e��X��s�e�G�g�04ӧ��|�N�Lzł���🻖UNJ�ہ�4��۞s ��~�YН���V�=ny��%����2���e7�:��o�Ria�dtD�Ԯ�!�C;���"��xB���)�u�)�Ҵ��Z7D<-�[s�Գ��������Y"D�1�p�5�u%�Ų
L���"�($�b��;�C�cA�AΥ�g�g�;ɵ\��޲�V�4]���!<gY�{-z��l0��d��7�ܕyZ@P�V��1����y���r��#�f����A�4��C����)�0�>��t{ђ�e
�s�'��ِ̾/?����s�
�6��Q��)�k'�!���o�n� ������ou͹���QT��k��Z�5Yy�#k�ZB��}�f#�ed)���҂�<�i�J��_���U�֒�D�Vo�ڋĤ ��R�_ݧI �,Y43W� C�Ԅ7đ�k�7���:��l�A��u���G%+8SY�dj"�_S1�Ɉ3�tb��ac�	�V��#����L/P����-[([�`�
�J��rJ�=mX���i���ʵ��Ύ���dxD������klv�'њ���\��1a�4��Փ'"$�d���h���߳�<_9���_�&d�������D��<KT�������c�m �H��w�a~���e�l*��q0���¦�I�tIE�A���\gC��Ӑ�K�J)�Ld���0�-��?ea���@	��|�3U�x��I�M"r�k�(�Cr�R�Č���x?=/zc�q���h.��a��t"��������P�o��u�� �#J<H[�C��
��&?� + ���P�`��y<p�d!����n������"��v�݇���P.2�tg�{Η����sإ��p�����K9�a��z9�*	Kg��9�.~7��O̗��(q� ���q�4�DХ�t�.��6����+�СC����NI/慢;�7"�6j?xJ4�$��Y#��ĺʯ��y>ށhZ�^��hɊ|�ѣ�Xk�lW��n�A��cG��������M5h�M���<Z$�RL�.�{wJ2�����)k���QN2��:=�����	��j5�5�ᫍܙlEͷT�W ��2�����(�_���ża1J���dTsF�(?@2��V���N13�Xe�tjP�����h6i��`�q5V�mG sPU��y�p5�M�v�����gA���L�����6�y�C"��z������%���;iYܷV��HV`�)��`7��r�gi�)xˍ`���(��8Q%m��J=&}}=i{P�m�K[l)V�,�-z�JS�͜[����/����E,�9V&j���2u�>��1�G?n{.�jj��H�K�=�]x���&#�e^*�8�8{�9�#�A�Z�dE�~�$꾇�q�p�x��7��NN�e_Im��$#�ټ�Ƈ���/2=�Yl�)�ؚ���9V���u h�a�fx�L��p3���6c]!������p��i(QC�>'�<�S�{���$��b�Poo��䓿����YwY6���T�O�#�sk���;��cY���qQ�G��8�ި �F��$3�XLL�� '�2�Y�$�n"b}��j�K��\~��r�q16��g�)�������HG�Ȉ�4s>r�>}��wǄæ�(&���'o:i+jqC��Jb��^������ħ��W�j�/����E:6K[M!�9 �-�"!ރ����C|:^��a���n�����:��?�j��ք�tr�/���l�ч$��aM�:�1���b���XU�/��! )*4�} �_��T�yp�Z?�A�wz�l���o�؀	�8c�nɱ����f�+��ӏ�]g 㟃[�@�.Y��s�P����az2N�;�w�+�c��rAqa
��a=�Q_�p㵝#?2�1h3�
^́zc$��He(+��tfJ%�mN�َ��rPs��hv�n�_��C�r��������t�/I���Y\�K!�e&��m3�(�t�c
������Nk�`x3h~�Ξ4O<����#���$�˖�*[j�0�� �YB����a�i��?�<�g��\:�7�c�-T
G�ֿ"	.�5��~��W<�:�RZ�5@���:��n	ʛ-��t���%��w�`����D���q���h>��$��%2��6�*��G�}��ɹI�8��I��|�m��{{e���þ�#~�(� �/��H�"Ԓe�2#��vj�A�rV�]&�7v|��;1r�O2w�
������C=Z���D�
:|���zʩՀo�����ˍ�9��	���j��ݩ��cgf1c�zht�
�ʈD�'Ez()"qN3��f���(�@Mt/LT
���
4����W�z�VT�#�P�qz��}9�p�ũYq�ī���ȡ�o���v�]=ߋ�`b�C&Pkc��Zt�VMA���q5�q�W��
Oԩ�fcpK�T���\c�l����i���s�!����a�e�[����&� "��UGԹ��u9X�b�P��uPa�Ćb��k�Ȉn�V����&���H�ٟ��u��ii<`�Q
0A�kE��x������,ǯRŤg���*Sj����O����89��D}�a(�Sf��:�8��:u�1�� Ċ �8��Xg�#��y�@�^�V��3d�����^.13�È���Ә�*�����\�$��U#}&���Z�J���K�Fo�K�������T,8�������Ecn(f�	��HL I=��ہ�xlbZ8�$��}3]�KhD�S_�4��~'���eƘ�:�R\��ɋ�=q��*.���}aӚ�
�;R��&>k��i�?vC��*��-�x�6��k@��A�F>���>��\4�ֱ�襎�/@͙瞳�*�-�]>��f氕�v�(�?�ya��L�z`��}�y�N��K���uO��2�ۚ�"����a���@eΘ�EϽ+�\�%���IL[�[I�;?�վ��?���Z�F��!��T9��}�k�VL��P4�ߛ
������������nj}�DՁ���������z/d��m�!^V+���߯,�;���'|��eb٦���=V�����Qӻ�Mjes��lb�cr&���GS�d�0�T�^sd��ɠ����Zlb�j3�ᷨA6#����2�9-u�Z��Mi� w��lV�|�o3��^� ����Ƚ������̕�Fd}V��^1bx�.w��6�j_��n1o�ȫ���ۣ>̀��&�rt�U#�u~�!r8�]��E�o�!��>|җ��1ڌ��l���C�#bW4F4X}[�R�^bS��:�<]d��t[s��#��V��d�������V��;R�h�SD4��2�c�O��(Q}ʧ�uPg,�d [�IH_�1���h��S��KE�i�]�{S��4љ�_N(�q�0u��?�I��YY{���Pn�?%z���)�TMR^���L��ö�qI!�u(C�zqe<��j�Sh�^=�w5�ϦIC<W�iIi�5֐Ў.�)����O�caX��|�����g�ղ�
�6l��뿺
�֛aTw��%�ց����-J���.&XC:}�4g#������y�Θ9�e�a��mW�
��G�7�-���އ�B�u��H}*u��7��Qf�bL��M8Z%>��L�m�͖2d( C�ii?���E���3����	��B_���
#!��+�=�x�YB���0�I��ab�ū���i:���ܹ�mkDO{&�]�����cҦ[u��ˤ��A��"�N��E���mwn���|IbZ�1sV媛�K*|���&Es����H$�&�2�7�ٹA�1%�;�&V�Kv
ص(��B��Ƽ��2���|�\��ŵs�W��X/�;�#��cd};X��l&�d�DU��UH��m����x��cꀷ����,�U@���m� �Ͷ��4��4I<ߚ؇�D+:��
̞[��/��x*��!4؜KZ?�U3����'�{l~]"�mj�^y����aG��6o^���.�/,ػ���8�1���R�Y�=i�ρ��ԗF~�㌈S?F���^��B4�[+�"�-��O!�fD�����	��=��*�U^���ܵoX��-)5�`�0B�L^H���^ �e��e��8����FrL3i%�_�p���w;�}6���ִ'�{��������a���vP4�ā����z�dgP���CT-�������\2�82 �������^/��ʰ*=�/(���T�z�,�V��<@<)>8ا���0�H8Ƨ��{r9�M1���&���2���2�.=8�>���l��X?w2�(�y���oӡ��/~y�=����,*��<�dR�Gy�䔝=}i�@�K�Kc�M�q�W��ʂ���D��V:0k�KHd,9!+�w ���?'�l�JNϹ+P����"�?d�r
�(��H�'{i�J�/D�Z�A��F��U��U)}�cك(`[��L�H���G�N��y��>�:�t�r5�mK>O(���A���Oj�;�����AX����p��}�7�-h�GU=8�_��l꒺B��mh}���Ln�Ӹ�53�}����uz���P�t����,��We�Zߨ޹�)�'�2l T|�y5�Ts������{�۽�F���֍%X��L�4�1��lP�n1�IE�\|uދZ)�b#���BV�眬�\̠֊��e��ݚ)���M��6��z�	D0����,G�A�t8�qz���e��Dy.�5�?�r��ڟ?� ��ا�����{�td@��9�j�V��*�&����-]1�a�o�f�P������K�j0�W~}]7���
�)Gk�����n����R�Qp���1>�Q3_G���;ͩ*
�	�~�M��3���L�ua�
��1:�m��H�ُF����x��	<�����*��R������}��+�v�%��yP�5y{p����T C�y�2�+F�L�*ko������^
N�F}(:n�rp��bY�S�xL�񪭏�Ҫ����m�@�qG�"����կ�����`=w�aJ/f�ih�����Q��/�k<Ji��oV������M�fs�D��ݏ~,q՟�]k�nT�1����j�̆G���7�X�xo!�����m`aGK3�y�v�����N�t6c�1��2Ƅu���Nu���FS��+�!�%�H��ꔸ�cEf3����8@L"w#}�<o���4�WX�$�����e��E������;t��q�P���4i�{�ᤐ�C�U��� ��uLe���\TKL����m��Z��{�|��SN�K��r��p�A���Ͷ�ZO�R*}�v���=;�u��{N��"�i411|�����ZPf��>l�80�Od�S�A�.cm��7���i���nW�1���ĹO�r�3:xَܝK&����x��8{v|�d��7��Xb!��\dT(K�,�֊��o6q��n�aк?�7�W��n�p`!W���-�k�S������Ŋk�${�^S�\�F�H��P�Ou�����kQ�#�m��a�6I'��^�rvp���0��)�Gn/e\1I�
��5�8��#T��g��x7W�6�M6�GTI�?$�.Zxd�_���N����I!|�nP��i�MJ>�yڡ~]:�A�3 ������[8�R�Gw��h�L8�} Y]��j���l�Ӻ��V��,�V������5�S�%���Ł�_ڟ^��vsJf�������ʉZ�g��|�·Z��w2�_���h�i3U��N�iǴv&���x�j�4���#���S87s���В#���7�����\$W�EP
Қk�m��g�uޅ��+�=�:��Ck>=U �K3��1�R򵗔�|Rh��N��F���"����IgB���Ux���Jw+���d��{��Oq����݊,{`-�W;� lQ��|f|mw�pp���`�ǝ�_*�\��0�S-��L�1j��1������3?{h�cRGv�-P�X&��㫩[x]C3i|�3�{:v�y��ޜ�>����F8���9ư�3v��2c(
��-�G߆ɜ�����'OVX��mR�n"is��-ܸL�G;����^?�@�1���E����|�M���7����K����&�si��������W�j'/b��ݲ�"�Jȹ�n���2������%h�]�.�X����N9J:׽� ���X���y�ؾǌ����*l��Jx�W'�!�`�nI�\6?�(-�P����Q�d#L�U��m��jR�#���}M�4.Y ��.�i5l�ա����Ɔ�՜���h�;�-[nr~�G0�>��PsF���!��Z��Ӆ���T2�A]�����*�j��ֿ	�b�o��3��to�8`@�d��[.D�Pi����4F���n���ޥf�3�1�&�դ�����AC���)��?��Ӵ#�z�`�W;��V}�P�9���F|�u%�ح���#�:�F��
�*�$ v�h;�y��I�x��w�2���3k�Z[��^ma�5;} ��f�"n�S�_}�>�[�)B�� ��'e��]��H��Plᲀ�J́�Nٷ?�kҙ=�q��<&"BCAT�,X�� �`��β �9��O0m/aah���!����T����a��d��qqF���=��_�\�H����������3lG~��Rj��.JPM���w.�0&��!�m2m�[�^%��/?yo>�,9E��Vb�U&�F�3�܍	��a�p���?��ŴR���
W<�����c(��*������|E���K�7%��J����I&�mZZ$M3�#2�b�s*q�S�N�dH=��g-��28tϓ�]�]=R�m�Ѱ���������iX�pU��y0�M�g���+ԃ�&�e�@�����?�ܳ�̟�C8�����b��A��j�MB�bb�U�{���A~��o�c@���7M�Q�!]eEJEc�S��'����U����=	-;Ә�n�l;"�Å����{@�k;,�5����$�vIc��7\Y���r����1Y�R��7�ьqg'�����0�L�%{�;|:1{�X�_w�p��c��2o�Ԩ���s�~K�+4\��N�`�������6me'�~@���;�������qi����f2~A��h�K҃Ig������Q��
�D�l���Ҿ����� %��k=��8�193J��4+=��B�/��Y"D��(W�Y��:X��4p�[���S��|!��6ձT�1��u�$����� ����.u���4X�q�kxŏ*�N�V�od-؀(�3�en���a"(t��|W�CE1�l����x��ß�g�����q���~�ox��#J��m�.��2yqmW{��'O	���vc�H�"n�>�����C81m#a�Uٍ'ԊI} ��Bj�s���43i�ӕ*���jwsD7�"�i��i�Rhp�����4��a�����O׵G�dc�L�M�<ѿ�p��<4���73d*�N�>D�g�*��R�h�3�o��C<�֘��тέ�)WoS}�ك5g3��&��I����[��~L�gw+�M��˩պv���\3��IL(����#���~I�΁���:ӾL�c�+Ș(t^�����S"����[�n
�E�^<��&��Y�@�	�2X+:� �}�d�DsC����1�N
x�%]�ͧ��?z<ȑ�����'������MF�� ݕ���ݮ�=���HjQ6�������5�z�A?4۩ǋ5�W-o�U=h���ʴ��M\�8�{�~&����@�k�}LF���,5F�#��tNX¸�M��-du�\yLՈ���<>oE���ͳv����>�`���M���x���$L+��^����/VR|��T���c6��݉q�m�ԃ榜tE>nl��� ԭ�G�3��m������T3 �{�*����gZ� �ޠ�]�J��m�HZ ��e���>v�j�{q��j�Y�.����T[IS�֪�k�};�_�B ���K~R��7Ym�zsOU���G�Lw���<���W!�B��j������k��.�a�t�|Bz��)���b�OH�^O���
H�J:�?�Sk��9&d�У�!��&��S�!P������q;�H�Cd���@[�����@�9�K�JH�f���\���Zy��v1�H��)�O��7���fCz�3#�\�he=��7��� J��%��������7�iŗ���2a2�@CN__Z�>:�����D��n�y 2���ziԅ��0�:��P�Ѭ@p� ����1�պ2Z}���>��X`3o��tn����Gj���^9���;�z� ��}C?\D����h��h�p�FO���u;����h J��S|\gk�U3�}��O�;�����w$�����3�� 8Á��e^��eg���+���)j�g�ط`7Uuh��2#�n��ŔK�נ=x�n;~)[7[�7����z<io9�5��`F����x�I��38�q�� dDA�bn*b�i|�D�Y�x�����v9��nvK)y\8�hY�.�q/�f���=@��w���Z�Y��
wW��X�L�#{xD �7F[��!j@��u燱�=?c��Zk�t����q��Y顫e';�ɧ;�Rᱫ^�Q�1�^�{`=��Х_�C0�����QXb��u3D\�ںK�1���a9�>(��;�p��.:��K�~����$��[�/z��dB
I�ܝ�8zp��5��cJ3MC��Խ�<b@��6�Y���b���L�S�
ICɂ�r$o��'���]����NFB�;�વeI��|�A���Q�q���<)1%�	�O�������n�s�]׀H.�&����A_��N� 9�	mQ�� Sd@td���i9Q����x�p{��o�a�#)*��2r�o���?�7���A�wCqK�v�^�I����)����GFY�='I����rU�\
�TT�Os��N򡘩DR�P�)˛y��_�7��&R��M\j7gDft{i�����g1
�I��"�S��(.���s #�Xo�	j�x�l�h�)����Q����)�Eo|&g�U"݅G��p�]��������`R����2d��R�����@F��*j�Q������+�q@�6ϱ��5�y
�*,�>�ؖ �@������YW�����X��9�h4�s!_��"@&Y�L6^�vye�(6��)�k���[;������H�R��ֶ�������u���)3DF?�TPM:��	I�����6�/'���"a��{��VCOb�=�5�_|f��*BS���L�����OU����� \`�.[���~a�rGV�*�%v.��6��}�L9���L%8��M��A�n��S�,z��9Z :lǊ%���J�ii2����dߏA�ݰ膬8����^��T��㐟�]��:����v��p^�m�+J��U�IN�s`M���fdY�If��_�a��zZL�!3��M� Ƥ�_����(+����0�sC@�+�U0V0�G�)ݞ?����p(4̷)�.;ht�S�����.[U+���69�#M��w(�6��ܭ�$E>߼��@�M�:۹����H���د�y���g�J"���f�������b���#�(T�1�+�6���$~>��XzO#����ۅ��(�2Vx��h��d� ����fy��yJ7�駺*������6�u�p��O��R̼��電�D>.��N"n�+�=���!漌�I�~E��e^)����)�����
�VC�X�
��}C����Κ�x��B�&&ID'x��v���蒵�ј��:�s	�3D�|��VL�'p��N�'�B9GR�ْ:}'S 'CP������8�p��Ao~�g��O� ��g1z�J�覈�#0�I�����F���>�k0]ѯ�P�T��%�3��Q<�cjb.<�@�z�W�|�m�t�z8-��������U�R�(c��&�5��;�����&C�����[�-�n�g�O���4i�H'BS�H�Ju�}�����r����l]�����C��z_���X���@H�@MM���o�n#[��\Bƛѷ�����s���b�I����;',kU�8��}�֏��G,p�s3Q�QG��&�M��`ڼH������|c��Q�0wa�TY�_ڇ+�oZ�J�����8�I�Q0��Wڗ��Xo'Vʪ �O�N���<L������F"g���9 m�^�I�3'�_�|��]��Kr�����"�D��L��l�+1A0�޷������Qӓ��<����Y>��ʮ��g��;A���z�+�`nte�{C&�w ���b�sHW=��-�f�=���>���rD���bԜ���G��&-���h3�J��H	�?��Z9���,�'���FN6�p[
A,)�Ŗ���2;�oI�:�:4/�GuW���+C�n���;�6AY5����-��^��(^
�XFǪ��=����cm3JU��@�Is�������e�,�p[ �����	LI��5g��Q��&��YZY�Aw9J����g�+�D|����*�UTy1���,�C��g��e�j����/�%6%��#�`�ݞ�\#����5��	�M�G����Eݗ�U��%�ӯ>���0��!0�cmX⤥��Z��:���@����q�#� �1*�'_:�4�rݧ�B�?B���?��z���t>����^�)�ϳ�(�X�����X򺠤�eM(����5w�+!q�S����ѩx�o�ϥ�����p��}�IZ���P�tl���	Ѽ��q
�9�]3}�^a
҈r��m�/��f��l�fTЖ��׾�|@';�+��(
B�ߴ��/{L(�s�l�^�5���_S3��<f�F'����Y��������Uf�hG��]�^\��vC�aYDb���݉�����KbS�%J�)6��D�>cc���C���^����Ӝ����U��{v?e��Ŭ��:y�}��L)x�as�{1M��(a#[L.T�5U�x��˽�E��P�l[�����ug��fR^a�ˮ	m��7�lhޅe�Q4)_�kϾA�µ]�R�}}�$���U�r�Y�;���«������f~q[_r�'��M�[I]���B�H2�Rj��
,ۊ}���>2���p?ȷ��3�ea(�&%�>C��']	VB�TWђ2��)a���,ȓ�ÉR�P⨣[|��qa�5s�8hH �C�x�����ɂ\|?|�If��CT�1n#݈�E�o~h����b��|r������&���yC�_쩱GF�$i��U����l6�s4A�dpO8�������)6Z���@W�y���%����/�����0����u�)�aR�?�:�HK�Dʘ�U?��(!nO��3󂟷�d��%���~Ǹ�,nO7����1nC)�� h�H��4�l~�i�d$���_���Q���{,���´d\p^�~�6����
y�RH��ۼ����.RR�D[��|�Ɇ`�,�/�WX���M�,�2T�H�kr��C��7�G@'?g1��ࢌ��f��Fb� @�@��׌C�X-'et�"�c��g�ボ���BG��CUS�qb�u�:�xI!�C:m��M��@s�$�j�X����G���q*6���n|dθJ�t2V�pб��Cd.J�ߪ��zHGd�N�ʻ�ٱ"]2f�8DÑ�F��Ku�L2 ��O)?2)���
�2�R�S�6���L�'����� /_��䤋c;>
�������xZ�>��}�F�T�x%�#��Jq�H-N�K>�*;����.���;�V/VĪlQ?�tu&����7B܊��E_8�0wI���I�����|X52��S/���9#� �Tl�a��N��<5���>�	�9�-�����	��/Fe�T�xx�թɜ���4��h�Y�V�ń�_��&>Z���2��O�5�e��� �$�T޺#R��~��c���@�ܓf���-+v�+����a/:�����D�����Jf�j����U�O��(u�bK�U�go�X,hل,?��7l��`����7>t:��l����#M���>�����-�3
ג�-	v��L�v�)9s�Z}�d���&����Z��D�/��5y�Nj�u���r)�1)���rn�����c�K�y�J�M�ȏ2���0{�>��7e���2CP�~Ϩ��k�Åc�+5�t�9I�rA�f�7���	W*vC���?*,�z�p)��cF�*��F�/���YӚ`�"��a��������K�9�����Y��Zi>M:kH0�k�w��"�����>�w���r�	���$���4���.W��*	N������vf��6�G����L������>���F�wF۱�r��᫢���jl�!d��^����g}4�� ���r�_�iR����eE��L����mx�v��^u����їm�~�k7˴Ɣ�4m��K������I��LW$4-]��@a�4�C(��]��8�9��|�PZ��ł�T*c�V@�W�Π�CU>,a��?��8:�*�,rɹ5Z�Ð�?���8L�ө�s=�Ԯ(Xj%��[D`Ϣ�
���`�4��F;<�a3��}9�3��>_e�,~(��.�H[�%@] �\������:�6֧�Q_�v+�[��j0F�HE����g��nk틶���Yy��A�'����qIݸ����Z]��n����9s8KD-a��<O��3��|ׂ�Ӑh�e�|fV��_N��|1d�G����
Dy܁[�'�uº��%����������c_��d���]^��2g��ꭤ�GJ�ʹ��^4k����d�P&�i�M�mA5���h6,@]d��4�أ��y)�s1G+��� �l1j��!���x�F$ a־����ھ�+Ae���SJ��t՟z@��m�o~� C2}ظ1iA���ɋ�*�|��:��tEw�Qݨ ���3�L�����0ȼi�B�c���D~�I���G�x�g3+V����a��o���Knh����@}n֒e3 d��@���e�O_�/���i_�x��s}����G�Ehs"����Q��1�Zt~ n�K�-�����^n�!�:k��6�_Έ#G�ټQ��`�k5�3����w�uU	ā<i�hA���iY�طQ��]���)Srڒ�jc��b�Z#Н̅���u=������=�7����t߂)O���d�F��Y����rL�	�ݴ�*+;\�pso�ul=po��"2m1�� ���
���Y�݈ ��gS��ɉ�S��F�9lZ��T! �eC\'B���ڪ1C�Յ��D�l��|_�!
ՙJS��b��='3�&���,-vW��գv�S�g!@�D	�A��!N��XȎHRO�ۛ��d�Z/l?a<��'/lTV}��M!�ΆZk�NN&�k�2|v��%F6u�8Fо��2�_�H`��ѨFz����b0�`���~(�Д��d@ؼ�2���C�M ��հ�{@=�k�9-�?q H�	������_ol_��BD/�y�:��{9)��ICwF�� j��3�F�P0!��v�-L'	"I���e2�/gB��a�2bp�luYf�a|-�%|�b�$� �B������P?���xM�P0k)2�d'!<�-�,O������(�g��#�W�M5�-�X���a����-�Zr�\eZAx��Pg��\ڱ���&��.���e���
0���SUA)�N�~���'")nʾ�!ԝ�>����02�s����)шZq�R��	Ѫb�w�RYɲ8�q�>~��w>o�o�Ha�ޞw؈*�s78XEv�g`�wCq:���~�}���l�둄D �k�]/w<RJ4� ��̇�1&!X�~�~+��bgg[$'2��{c��E �={>�u���J|��m|�rB�y�f���WԠ��!����GX֚��W�v�g�G����d��(B"����$�/�0b#AO�%D��߉�s��O ���ma��`|7T���l.�Զ=����(TC���C��>XЭ��Y���E����~f�dG?R�JZ�~��L)��n�Y�Q�} O2��3 �T���T��5�^�M	H�9���dy�᏾��ϙq���ŏOO��*��}զb �@�����@��lm��!E_����U���?��M�,I>x��P��8j}�I��.����-��!C+x��]���Y������eBOM�A)s����5ؠL4z,w��.U����}�^`�TkQ6��M���[4��5��ɸO^>yMs�� �L�ۛ�����lϫqS)�bB�(y�q ��딗{��yڌ5�#=�K?���HʍIa�xFL�o�(w����/�����(���U-�wVb�7�a/+1��vd��g�K0��R��$��[zj&��X��1J�S޶��k5�ձS9Hr%x����CڔN�!�@
Ҡ����Y��A���}ᓶ)�-�����}��6C,�`��O��l�6���75?�ڲ���'�E=��0R�T�UF*�+8�#ނ]�3�`!�U�L��TÃ���	�K+w3���s�њ�ֈ��"�c1�����
�����'���a0�1T\Z�o�h���.��93�U��}���s>�9�Ǝ�2:`�,�N(Ϭ����4`�*g-�T*��j���g5 �3�>8f#�+( �����^�͝(8�� i�!��&��R�s��\�n~9�腠�x>�e�f�O$l�Nx� O��~/mS���# >�#����9Yp����Գ'qQ	�O�����?R.�ڏMn���J���Z:Css�c�w�q���jl�%���SU�mF��CLԬ��I>�K�q���	�2�l?ӯ"A����co��+���A�����tҁ-U���?k��\E_R	��XG;Λ�Z�D���:v%8�w��r{2-n�]g�0��� �L*���eQ"�=?��޲(�o��� 0|RDb�L�b�mKr�m:<P��j�2���r:�=�D*�#p��8��C0�vYc ��F&8W1=w����w��E���2U��q���G���e�$D���Z1��3
���I��̐q�j�jUɠP �A3����T��T�Z�5e�(G�2p����'�Wn_E�p��&ܦ.�gA`/J��;�����.e<����1y�Z����^6�|�hh�"m�1\dd+����<~��%
:�`)�D�;!�k��"�ڪ�Y��5ۨk�,�*������9�C�2�����g@����|���5-������n}q"ϐ�%tA[.�3k�SU�:7ڻ�PR#���HF�	u�����<�}��l	1�t�EO���/�q���?��?���kO�Y�iQE�sW��a�+�[G�t1F��e����[�=2\eZ�r;�7�=Yw(= CʇRܢ�E��F�K��\��B,^�׌Cđ	z���ߔ�C�'�,��=�� lr}�]���3�=qu���a�ľ�������#R����D��	}
!�<��� ���r���F��7��J\�b�n��e銄:��¢7#/��'�wK1��:L���1�?�;�<��<p$��n9�#�k�q��{�&�>[�0�{�Q&�2����u-x+9��!�A��Z:i���4���~$xI����jPYĜf/ǎ�u��h�R�*���~N���u8�;��h_�e3F��"�E�&s���=���}�.�تm� =�����Ձ�;m 2���K���8��,$��9���q��^%�\���uH����uvؐ풒�=�o����v6�.�+z��3_��}�[�����bw�@�NlW��������U�L�K�F���潆����~~���*�5f*��Xo�����ia�l�hpuq�(lo���a�H,;�3�L�異�J(ZH��sZ��5e�i{d�ZM��.=�A�l����h�������xٻ�X�f�h_4�'���Y�^�{
u!��	uPb�:jG?��)����nr����������5��_&����Q-fe��x8�Ѹb+��bފK,}tf��]��W��l�~���}�6i{��Z��$yS�qM���r�.Ms�eLP�������r@[�
O�Q\��8���R93Ђc�B $O�|�^~�#��s);�	 ��^C TC.+�A������P5�,ɼk���M
�P�%��n�6�9e,3N�h��G�}��ytt:��T�w�g@���bJ�!���.'�\xV��z�5[
�n[���/d���g�"��I�Ʌ�XoЈ���v�&�|H�r�~��RLh&p����	'�$�NxL�G�GD��5��C/.�R��L3��.D�\~��d���rB*�[|(Y�
�?��9	��A瘱�=��0`��\�#��=>�R�d;�a�����[}�.��^Z�X��`����r�-{|DM����"��ޞ&JL�2�V�uh��	"���~�^�Y��Pr�L�ߪ�j֮T�ױ`?������0�1�����V�w�\Q�p��Þ!r����2�cT�*FH~��vT��j��x��a�t{��6��d�0��ޕLX���<�)-����\&2�A��e�*7��D��!�@�R��-��;��᧨U>]7fx����~/DSڰ�	�m�.t�'{��0Ϭ� ɲ�*S3�j�Z���{�1P���K�����(����u!��gF<�g���lg�f? �����`���%0�Yq�
���*����&/�&�݇�oJ��;����]�<0��O�N\�9dȬ��:B4�%���ش���*p��3�!��v��U���'m���׿��
˖m��i8k2A*�V�Q�����@l�?S@�����
���3���G٣�cS�V9L4ȅ#ڜ�u$Ay`~G�����.��f�MxH�T�+zy������0AI��-�}X��-&͂��{V�ܩYjĢܙ�!�ڹ�Qt�~g|i��
~��E�_;MX0?��'%iE"���ީ�~�Ks�ߒ�(�o$��t��m\�n<A\�:�n`�y�J��4���2DbG? ͫ�Ѩ���-��XYZ��9g�
d8� '[ 2#▞O5�D�P���H!��z�_����.!yŉ���Z]P��t�����}:;R*}0���*�^]T?1p�:�z>�4�VT����v�r?C�ul�{e�kd���KB-���I����h�/�/�_����o����s�Hef	K���I2�w��R-@Do����=H�P�k;���d��p�
��$ O@�C�n��kV����z�;'����(�|ku��C���n��,+2���²���o�W���g�l������<����T���P�Sd>a���7����i��
�y���b��*1��/�+��R�C�p�L�N�<9v� w���5)fc	��I������J1ǩS�lx�H4��f�Y"F\�P�l2�@!8�����y.�0��??`�mf uC-7u�Ť�'�u7���h�� �`g���S�5�z��F�����z}�՝`};4��ຳQ�"�RHC��A��x����%_��ɝ�m��ifd�;wdw���
A Ey}�c&��E��B���D	������ݹC�,�F�$����(B��w<��9���0H���l������To	<X')�qpm�忐0^�ً��;$��/��Ql����4M�)6�Zs6
Ef�U��fW��+U����-۽>sp���b�؜��H��c��pO ���B�}�
���"���Gx���M�}�&��k�7<�\/�P�%�Zd������_E��aQ���\�I�K|e+І���D�V�]ڨjt��N(��{��PZg"����8X�Pv�^�,����1K���X�\)q4�qu���8)0i��7�̎�;�m;�Qل�,0�&����{<��#�&��'~�%_̈��R#d`��Xi{*��kmq7�z1M �TfD��ن(���Τz���Ǒ�B�����Ľ�8F��7�Q� Q8c^�"�"C�wy/SjDGBn��'�.������U�h���ra�y�T�*���&;f��0ST+��h����2/AX������C'�|�>}�J?	�e�!V�x��C�\�]������> h�؅E�s!eۄs��&�t���l�jOFh)�#�EO���U�mV�w���w��� A��9�
�מ�`8Q��\��~�X=�b��Q�l7w�M��mL���������������m���7���+r]������e�_ZY�&�f8�
R�p|
l6=��+���gqo�7Ƒ� ������Rj�6 �ϟ��je��CH>��L:S�#^��"�ڧ�Eu"�4=�@l7��WFw cG�=y�y3�Ă��c������9>���qwp��D1u�-[�E#�"�㳚:�B�����ً�"�k���$��M�](XM<��AJZy�@P�$�]�"ee�OSk*Y�{<�?|	/��rp<�6�k�J����P{��R�Xf�§4yYX�C��T�ۚ��]�UP{��J/�m�_�	C[��˰�h�U���,��B�sO�h1������:ZA���(��i����%%@a�q�o�s ?׍������Dp;�,ҽ��u
f��/7 �����c���.1ς,]ܸ��#Q$�����-��!������y�oC��PA88`ё�VU$��9&Tp	�@(hs�_!1����^B��y��|���C|�^��Ub�)ezy��?/U�S~KI���8�{$0"�jY�������[a%&�on+���������\UJ��6ӓ�~/�~YEěS\�Q"��y�Id8h,������+T����zFm(׾��sP�?��LWu�h3i8p�F���Y���'��'�S�I���������M�y�ouV�����wWx���7�ǅ@96�!�h��]0	�zw�,	�E��ɓ�j�7DgЎ�S��5.��-�1�ɇ>��J���[9:s[=Bs*X@��%h��� ��-.T1YX1q�cC���Nih�&b�^ۘ=���
��w�
x'�q'��N��3��k-	�U���Ÿ8u�ҁ�H[�Ȕ��LAN5^��̄Y�ۯVt��',�:Z� �I)U���t<\���!��3�ĺ>��#�y由��i-7iw]q�G����5���Yu�)w0oڀ�ҧ�(���;�m���.�;ڌR�"�:*z|2ї�t�L�sb�{q]�z����� ft��Q���0{=�%K�B��.ܕ��6 
�h��5r�������S��H N(��Oy1�� ��lS>���(��6�VtUE���EM��i�ݺF>�ik��z�M�q�rwZq�꭬E)r�Рι���i��w�ҁ�7��\���D����$(,%��׌�2�� ��/�Y3�V���	'lS��f�$����`�x���b��~��)<��sQ6�<�������>�c-D�+<��cϳQj�w��;��Ε��7c��Nƃ2ԝ�t��υ4버�n�>:LG��ΰ��O�P�E[���G�c$!�4quv �y�qXmm�~�~�D]l2��s�P ��o	���zo�B������ۘ�!zQ�u�\�|�v����Җ"�O9+��Χ!�BG�jM�R�K�v�M��|��"q��|\��
'��(t� V+ـ���ܑ>��e�/'��'��^q	�2�ǜ�����bM+��캱�a7�_ >��nc�'���.<��N]�@�TS?��ɦ >��z�����\�f��^M=�ؔ�=���4�)2/jV�v Ɏ�}!F� �m,��aɩ�4�+B� O�쭗Ƹ}���'ױ�⍤��C)B�V\{�S��~ª���N�5W`��a�K�Xv���e���2%�	B��ɂڒ�k`��-�{��(ED�>��cE)e��/͙��|%����|m� S>�z��][�s�'
�[��4ㄿٯD��j���t34s�*Ͷ�ӑQc8u�x��S���i��mE'Y��x�(�=&�L���ˀ��F��3��9�U0�~ԋ��;�gi'b���/ra�w�j�m��Vו�Kb�L4��G���7D7n��F�n�%Q�a��;��\�Meѳ��_�������j�$Dݕ�9.�ȇyc�=��j����%)R݆&{:�6)��s/f8�~4#�O���~5ǹ�c ��v��::����	) 8����۲C+|,&����M�W>bu�W�{&�5�C��$��9Ng�_��!$�x[G�b��R1�Bo��+�����M��>�u�6l�$ɒ�aS�{��s��s�]P�����$֘�bG):A��v��Id3��8����c���e�7)ל/�c��p�v������|��c��i�U8���2r��b8z"��C�����\uB�[ЂSm؆�N�k�mqs2���/^5[U(�XLL!�(o�.�5
�Pi~��w�.9�*��6�\^������Gk��h>��$��=�,WC|�'*IL�Y�/�+'��B�K��]8!�4����W�M�zx��g��i�����d� ޹�z��~�]�#ۏ��S�����ܻ_r@� �O���!��*>�yqw����p��f��x�ԧ#�	 �U�l۔J2�sN�i�X���&���bn*�}��.�i�u
Ը�����x
=��3��^�\T��yd�o)�\��! �R���z=�ǘ�~���pR�=�����Ov'��0�q�`A��i���$�n�Y��0V���|�y$�'�����Y����2��a�H6���)����{���w$���؊Zf�<,
d�a>�Eȶ)��,�רJ�k�]꜃GR�-_­�`O���W=�g.NՓ�n�aa���D.�[����d��O.i�.���A��e���2 v�!��ڵ$$�v���Ȯ��t������G�O�����@�s:��E�p�N�����u�R[��wUoa��&69A-��|%���L�t�wU1��]�u+��݌e�h>)ۏab�c�2��ި�׻Z=�a�\DH��Z\eJ�Ş�֎��S�	�AZ'#����ː�#MH�
�[���͹�D	r߬�sC�p�O+���>���**^�q���љ6����j6M%h@郹��I�ۯWPh�0���I�"盾�4���_�F�l1�vz��'��R�>f�D�	�{����,d�أ��#����MKe��G��-�ټ��:�P7X�/���?�-��J��/<�;����2Jz�&\
�D����-��s��i����b3H{_�����rN 5���)�XFC�>P�.�U��m6a�m�R��ƫ�3��`�E��.�j8N�,�S�n�3�ڣ|�1�Ei@�𿗴hn�wu>�]��E��=�Y�Lp�%��`{H+���&eds#EYp ��#ߞ>A��h�4p�p��R���Np�_Y�1e���K�cG��e�"��i�-zF���7�&-=��̒��=�T}�i�/���&��z��� W'���م�F�E7a��.s}2-GC�Q��ͧ?�U@�6���G���;�K��esdD"4bP���5���W7��#)�:%0���Q�U���F~��.����6R��;&���<iB�1��Ϝ:��r��Y����w�z����#�䡆n��x��<:6��5����2J~�C0������Q�
�9(�H.��q�_~/rύ0�x�	R�ޚ�/,�NP��C+��e��S�Em����88W��d�%Tk����4E�&:�G�L(.}�T;��tޟ��2�=�V&�fh]��(R("���'�R,s��������E�&: R՟[�؛�*�줊D�� sk];���؆ȩ���Y�e'r)0��@���������2��^'B�Tf�:l�]ռ�$����.Gx�@��M��\	���F�XYAװ/�X�1��ѱ��:�4�iG�E�Ob���Ƒ$��Z֤�!��O�@Ģ~!�a��+�	D��fL2�����I��ؙtnvtX�9;+r�/�c�5�b�એW�&o?"7��g�
����� �k�v�V����3�S"&,ZΎ� ,��&L�������d*N5�a,VjέY�].`� 9ٳ@:�ZjB���,��ǸjK��N�y)@�J%�k���Ϻ�5?���#�����c�����=�x:�%��~2����L�o�y	<n�8��Ѥ�xt[���DLGzA�Av�d�����LɅǚ�D*w�AM*���|��
���鲆5��da�!�@Ѹ��J���/z �q�t�wC`��������\��R��4`��ڌ-�8h��^#��Q(��;^����a��TY���\_<�)���Ɲ��F��fV�J�V������c� 8�w��{MB8�~s)m��.��%vT�P��;z[����֞�7��U;׬˟6�t_��~F���҈t���7%���R\����k~���!�/���oi�ϸ�o����0Y�$o F����H�vfσ�a ���b��C|E(Q�~����:R'n���P�wK��T�s=�ɞf	�	��v�+s���e�nQ��T������T�dͽه}�ml%ᑁ1D�sb��K*�{�����[�����B�}���-��<"��1	����yʾN	q�f|�f�iSB��kʁ�� � �^p����4и�ޠ���ب�<C8Iny<���߼/֙�H���yx�4f�D�G��&M�r��{�ݰ�:7�����w��ʆ���k�j�m|o)d�y�i�X$�~L獔�VVf�.����4�>�n���TE�[�n-@��Loo�3-��C)%D���T_�:�lK1b2~J�y�%�:��¨�ԅ2�>�/V���	�X3�4.�xFQQ~�����Orp㿽�:�*y��t �9�Ons	�T�I��/�d� sp �A6cfl^gz�V������J����~��K��b��^g��|)����ъ�	g���b�Q���ע���f�V8�n�3Kc�,� o�UbJ�N��Y���?\I�J��6S,��B@x���S�m1�0')Vv�����M��� JM�^�us��hZ��G����N�
�*��}�/��:i~q�A{x�y���]�\E�m�veA���	jh?H�%�;0eQL h� ��~�XB����RB��������ɕ����X����ÎG��g�S�uȳ�b�z9��&˔Y�Ob�L�#2���>�ڵ^�1�Ή���T�B������TF}�z1��vRV7�{�h�Ay�5�ƇB����`+�O���ʀ�bs�t�T������6��$�Άy�4c�_N�7�7b�5RYed�Dr���"(9�ZԊ����L}$�isEm���������VȪ��J�Y7��fܜ"��ڕU�������s�!��ć��%�B)�P_&��Օ)�w�ƖI��ш�v���o��ִp�R\���V�_nU��1v����S��c*[�7�����0�L�W"��)���lIw��{�O��l{�ݾH��	�\��4�6���+�U��r����>]EC��^�X�PJ$�(
��j=dі �z��Y�Z��8=������f�?���R"C��Vg�^�qD��#�#�D���6�<����f=+Ȼ�,�@M[���E' "T��G��ۉ�;+�9�h\�����U��k���R�����d�1Ş�_�F��g�2�&<4���P
�R�*K���V@B��p���e?K�tV:�x�H��_'P'V(9�yu�}+� ��|ۭt�B�[	�~Fe	G\bvx$D��5f����q���^���hG�'��߰=(������
�s���<�	@�E�/�r�KI�9��%hWz�?��]-����#M�ߗ:O�3)��\� q��߃m,����*R R�|�j�]�R��c�M:��j�$�NOSE&j�Lx˒��쪠m(���M�w�)A���j�ڝE�ж�� kf��x�J�ZFR�d�9����rVl�c^�r�wP |H^F�ͦ|�m������p{ڷ�V�'��Z¼�h�`a<"�1QVT#�~+z���>�1���W���Id�8[��Ǳ�F7M\�H���EG�93v��T6/aД��mn["5,Ƣy?<�6��v<M�9��Q�bl�&��K����>�ޝjŬ� �0��X�@�,v'Z����r�n�bY�c��!�S��.s���Kc�o4`Y��}����h�?��~Q�͚X�@= {�p����
ϭU%H�]g$T�2eȉ�.L�z_k�)H��O��nJ3��b�-M�@fX�����M�%C�vPهk�����<�1�pԀ1�WL��T���L�w*�8����[X�S%�ؓ0�eyDu!t�zk�m^����]��y���f��D��!�D�����66"�(��MZ��8�����s=gw����b{ǀ0m0 $��w9F��z�d�s���m$��߫h;QL�z�u��5"Ǎ/j����ɯ��J��ȁ�ґ'�_�:��<�k��S2��^h<��kh�~��d��c�<
��݉�$�5P�\7�l�1��
�k��s�a�-L�Ƅ(���S�H6�#t3o �����Vyo�dp��$�z69t�?�|�p=��f`�d������$	Q�
X�3�
C zN�wL$��zD��3H��+��r>���QSV�?�*L���f	���u/Y�
�ύ��o|[����0����/� ���ٿ6
���Eᅃ���5[�v�_3���\������1��R�U@�l��Hc��،CKW��X��Olf�Ek�)�
1V��.pC��CC�~�o%T���8W"��P����R�7�Ψ�9^���'t�1����ɗ����_wӒ���n��h�/� �9�ԝ���h���Y���]#t��.ܷz�e�M�vf�4^���sE�����;��L]f��<��g)=A>�[�fS�E��H-Ƌz�VKWH£n;�OE�9/�q�ث�^ �U�!^i	/K���`9�EޤlScjiIwڸ�dj>�9�k=��-`/����oU�"@��f�1Z����O���RՈh���}a��u��S��Mm_Q,_�E���%9���:��ǵ���hf(�n��,!/��l�=����(R�f�!��_R��A*�t2v� �#j�t4h*�Td<��Ğcr������*��-}V�z�0�"�Q��P�_����b�l��r.Rg{�-���h��2�W��Y��ø�=�����P]� �&������϶ٮ�;�xk��{���6Y�;�U�>) �:���O����)�x�3?:Tz����c�1z�i
e��M���ug)� U�t;�<�[h�����N9� ̈�G��N��Q~y����A�$��W�H�,%(Jr�|,�<n�0^��j4R�ap'�$x[�·8� �-*�D��&T!ݹWxo��2*X��2���Ʈv%�|��ֻ0V�(�S�&-�)H��BR�4��X�Wu���,V5��kPdD��3k6�6���?����b����{ܔ$й�\���z� p7[�]b�Itr$��{��g�u/���I��Z[E���ח &��|�)�цYs'|�aEZK'�C3�JU3��qb���\U)��M����xu������]Ɣ{96+����jtJ�".w�dt�B�~�\9��̑�[?���È�u}������c	���<�[r|�j���|���w���sHwp&��ЧiS�%Et��� �j���#4F�f9�}h_�K�[���}�����8��[1�0|Y$4��v����,ũ�4�|6��}�������P�D'�z���K�`(\f��O|��hQ+��)��aL��i�4�r��q�U��a�'K��h����0�w�e�m|�����#7pr�o}�K���K	H!�-A�,Ӻ����r�<wy���T����t��;,cVx���(/��f��B�����ت�K��g�^)���g(SΎ�����78e�>�w/�D��g��%/L#s0P�)@���yP������M���B8䲏,/�oC�Y���LA#�(�_��|�X� 	�7�
PiL�+T�5�����dK��	%s�b�^���GU�Y��`{��=O1�I��n]K=w�������zku_*�3�Ƶj@��e6{�LF��%^wa�`�	��vN��J&r ܖ��]%�a�[jpF��?�%}���`]9H�����\�u�6�0�m�U��xٰ��Ȏr�ʹ����w�9��'|q��,a�Q"���n����E�W�|H�7k�Q:���fP���
�60\��i$�	}bT9ZwV�M8�1ӂ>�EF�-N��QB�6~j"�fY�����Z����J5�c_m7�i����5A��p�郎��[����W7�L�A���8w�7��E�~O�[��-0+�"�t�*�GC.�����2>R�l�>'y��~�U�ax����S:�u0dw>3WI�z<��� F*��1��F��B�v��H�ªz��k��g+�3�����u��l!��?���.Q+��z�^�}?7����v��$O{&r��hF�AƑ�VB7[f�@�`���9�l/��RL]�J>%6�iJT�5H�����}��8�ʠ����h��@ bf������Kم.N��v����Sų�Z�h߭�k���Ҷ����^oL*v/Fp<Ic0�b��ɚk�Cs��{bhK�t"?�E�_b�98Z���?�J~,M8�$`\J��}n�������FD7f�=��k�ȷ����Y�;�V�T�p����0�#Cs�)��o�-\���o�^���/L��B�`.ʣ�{��+�i����B�U	C8�=z�+�VB�o��&�[+�цm�9��1�v�����{���3�g�b|�5ʭ2���
# ��c��<�����D��`���ɘq��,���D�	�!��K.9>][�Gk2:u�Ŝ���=��[��
�ܯ��L�+�7թB#�c���L�R�h������wy5S�KI��QU�b��}][j
w�'ܧK�aF=�aҨ�_��e��C�,�z�E�� /QU=���'^ȇl�H�䣅R�P�(ܣ�o�;Y���@v
:<6�7�K�u��2�}�/	���mTR��l���{��>ɗ�7�B`��Dm�p ��d��U��D�Ȟm�E0ɽ���ؕ�#�u�(a�.��zA{�_|�R��J���1z?�5N���}���%x1�ڝ#�b|� �v�P<��"��GIKވ5�9��MƢ{�	2Km��� ��Z,BV�KL"��^��}��OB�C�F}��g�C�U���*���l�-zC����'�\���+�_b�8"̋A�Nr�5���E���5��n��U���:�JiK�n��3v�1�e8�6L���� x|�w��w˰�����։V�u6����@�OʫX9G	@jSf�H=��W�uF���#� �Yx��J����{�[���/�`z�l��ݺ���\+7Ml��s�!M*V���emC*�U
e�&��^!�)G�kݪ�Y�N��8�@�M��6^Z�������Ax�e׺�ӓ�/R��_}0y����a/	Z�w O#�)Q��{��5��BFՒa`E�Ѣ)���K̎nI��_�s���v��)�J�xn�9-oͭ=y���GX|���g�Bn��S�;2�\��bF7t}"ݩ+/J1c�sSܯ�-�<�&C������4����p�I[�R&	uV�aJ� �nb+��n<��~�y�-S�!.�&cq�7ue�V2r����ÎwRë�ꀀ ��>�#£�i�t�K�a/@;�%͓:���{3�k�R�k+%��!/$����w���4���w��#�9Q	��������T���y?�QW<�J���W�j�	�g��r�)���5[��CŮD}�RB�m%&uBY�������G�<`����1���+���͟�S?�2��7�t�s�m���ҽr��_V�����쐭����k0���{�Z���h2_Z!<�"�����Q(���4#6e���~�T�0{��h��p�7R<��v {YWl��:l�W�:�.�(��8+�4�;����P!�x苷.�,�N���N��a[�
Gb�M��L�/t��M�Z����NSܥuk�ٳM_�))�P���x1fo9׿ң@R�~��ۅ/I����t��*bDj<��~�Y�j+��(V�-w��{�����X/�����<�e�ZZ�h/��b]H	%/�p5A�����@��Z�HT�@�������f2���'9�]*C�	��6ʄzD)	��ى�	iǒV��!h��fxx(�M�p�H�Q�����>E������<��i#ϴ\G��:�>�gS��*(�C_rp�|�`l��% ('��LD��������=qqЅ�r]#Նa���i���ܔ���?1*�Jj�����Cb�S������2�.v�EүsrcQR�Gq�AJ�����Abac�ҫߢ��چ�G�{1fb�19鸰�����)v��O�1_��g��݄�#�B����
�1��C�K$(R�����5���u���W���ӡ!QR�ȳ����a��cv�i�F�t���׷�RW�o��a��tB�3�Q �U5z'{����O��Ǩ,5���ˀ}���$���.����c�y�!����`��,.�K� `T�Md�J>,�5��PP��]�3��H�������Ҙ	�4��/����_YlC������&ꊌ�5��9�����i�͊
0������;�8��ʇ^8����'��M�L�>�~�n	Kj��W�[��a����Ll�F0�����E���#�rtcY�݁��*P�M&N�;E�M�Uzl�8�a��b���ųy7��h�+fq�������>�uCO�K��]��"�p�^�o�UK!b�ꍺ.^�������f�*�� ������ߧ�M��.@{�ᕨ��w}+�� b��m�������u��mb(8	���k�:#��DMMaW�e��j���)����þ����	��
~��,Ee���-�z��w�)�������vo����<����y<r*�ڤR���HKG�lUf�?�����42�q�P�Vw���g�:���>��ܑ�n�uk�\ѻ����X��4���䪺a���/?ч��y�\ѽ�w��2��fG����6�jz���0�uۅby�����R�.�7�Z%+!��Q	���eV��į������
#5��{J��i����J�#K��N�����{�d�/�� �S5nV�!��pm�18���G��o|����d�����H��B*�6���FfB�t����'�1?.�HK�9�hj�ez�0��\}��b�3�rP�`2�������[ؾ$/�ؙ�?ܱ,j9�����/����o�ǫ��E���l��u�h��	i|2��E�F��Dn�&���ܐ�t��p�>l�4���KLp�����q$��k�!�A߂�����XT������6�to�� ��!{��\O�5Ȟ`��fO�jʃ{9ʺ���ݝ����؋����iŕ�J��ɊSb�4�
�����P�n���W�k��367{��� �ڪ�Ԡ���Č�w�*q�\��
4 �
�"�C>:�����ʝN_z+�Tgy��/Db���4o:Bj������N�g�ٌ����T�G��\}nZ�����{�Q(�������%Q��!T[��v�.9C��5�r��Uk��+e;���ͫג՘7Sn~��Rn�w��-G�vH�!U�7)a}��&���s�m\mii�pa�W2k������oF�`.'��䇙����B�9�I��>�*bH�p0��veo���l�L�f�w��U}f`���\�=~:��t.��3r�/&x�,F�->�u���4å��؍g�&!��rw�ɦ�\L��l1Lf;6���z�����°�����Mu�
58��)(]��; ����(Fo�%`W/x���"����;�a6q��T��ۻAea( ͅx#���p����-��⾕ �P/���O��y@��w�/�'ٻ�t����"	�+�t�v��;���z+dQW��x�J~.0�s��XѼ��)�$EW6��)}�ֈ�.FA�n�-ɱ��S�q�5A��K�j��*�ᕁڍ=�Cԏ)�*k��CSeO����y*��ϋ��O�����*���n������>�At�������+I���.���Gਆԝ��P�&J�
��i̠6?r���c0Mgǵ�CX������d_e���<�,��X�}�� nKA��{T�����m��N�M�
$���V���5y>�ʄZ��5 �]�c	 �نy����\Nn�j��܂�ޕ���-n�!{VAl"qx��{A�z	�����Z�&����C�tu�w��`�.C!ΪSg,�0�,�%&�59�q'>M�oϼW���}l6p���"Q������/��T��U�T�a{@9u
lR~��X�&9 �h�t�V��c���PB'�Խ=sj�����qP�����%��\�%��fS�Ht��U����O�\Z �D��c ���A�Pk��-�
�A��{B���q�f�v�"�������g�c�%6�C������xRă%��Ƭ>��|:2�Q�/�Q�qB��ƫ���6Ga�t`�ݺ�BV|�z���y��>7�����g�
,��?�Z�3w��c?�M����q��tԶ�|��\��z�h��ٺ�Qcg�����P,|�E������_�Vɿ�&��z�ۂwW�%̱9�G�yqV&�L�D=E&��TZt|�D�ճ�c.�- a��	�]�2�F����8���`]��ZlYP�=H�e�a|Al�0?O�&�U�=�`�k�C�w���m�W����ԺfyK��n�*�Y/����P S�ѓ@;0uy���T;,Y�I��m���C�+V�ϛ�٦ �����MX!=�uӄ�p5c�eL�=M���ўZ�d��䖦-������b���h��C+H>\��.�?{�o��ylq���A:Ϫ��"k4�pd�@^(J,u�/e<7o��S����E�Z��jH�'+��+�IKD=��Z��\�X����Ʊ���� ?�����cԯ���)��as���S�.�W�5\#��ִ� J!�5��i�0�,0�!���>����
��!,s����
VdɆ��������2nmW�v��~T�H\����|�ܡZhGk�I����'��nN�P�1.�vGڠ�V�p���uF��e���Q�6�@�E�p��x��A%>e�n�LR�m!���yz��M�8$�0�Waz1&ӖKPR�YPpH\Ѵe��+��G����?��� ��VE܅��{e�-�����&����X�L��`dt����~�v��h�c�����o(�Af0���A4H�^b�Q�D �Uy�u���6aH?e�|w�dU��GW `�g���~����B���K�$���j55�͐ᠵr�W���x8U�����pa��K5��������;�PP5�/}	}q��_�r�FG���p?���k���n�'�����5p0�C�(ߧ �#T�L�o���>��A�lf!��/G�!�H9�'-�}��B�Ď���TZ5ը6^�ǥ�ڽVܻ���ʒsd��"���,�n�M�<A��*1|3��O��r�X_�ƾ!ma �:eK����4���'2�&����{�[�˓�u��r�T4>g��y�j����?q�f7T�i�0���$D^�yD��0��dՌ5;��)�K��Q�<Zڍ��aV�U�Aܖl�}������
���HU���>;�'Z���r�	�=���e�rN�;�1�X3`5-����gJ:B���"���p 2ܲ*��&`�1M�/d|�6���X����Z<���`�c }��{�-�&�e7Y�4�E�"F�� N�d��r97�;�	�̰��%�f�;!wA�0���k�'2؝y��i��NJ�p�F�d�Ő�8eg��t������W�����u�r�%�$$�i��]���	+v�ף*Q�h(e��)�{��:w^b�l������Օ5k�a_���#���Y����>����|�W-�_�mP�0VK�#�� �����
�\�m���)�'D�XV?�����u��捂�7�f9X�B)v��ih����	/k����Ϣ��
�/��h.�	7;
����Cy���uNfd�ڽ���܃Y?x������G�!-�'љ�.sO�c�\��T��r���'�h�i`�u�������?l��-�4%7�jOk�!E;/]�zVf�R��$�<�� �Us�)v\����f�)�8��El�1B ���� ����7�`H}��H��:�F%��=~T��ڶÇ�p+%����Iu��/�wA�U�,*Bձb��34��j&��9X՘��<d��4���U���`�1�,Q6Ae:}:e1(2�捒B?颐���\�c|���I�����;uѰe>{���F�|��R�4��>�K�[n����'����8�H��F�fY}W0�J�q.�+�'��ڮ;b!�{����ϕ�ܳ 6oa<�Y�7�<�y�Jh�Ӟ�/�ݡSO�b`���������x`�/	�0��~Y�s%,����_�1=�Gڔ��!���J�^.
���J��<���E"q��t܁-�n;X
og4�	'DB�~Ci��@Zi3�����!O�%�Gi��h��ls�a=s���su̓�Ae��^��1���ò{Q�B+4{:d$5.O�>�]?����=��<���Q�.����*5ī���*��j8�ąl^�E-��|��^`�f�!.O��Sp�-�+R-5�Z0�K�hڳ�E"A��Yt�cf%}���bI�	��窇��!�\�:��3�hN��8&�Ue��V��ՙ5����/�.�8����[���%Dn$��lm1he�_Ne~�m��	�e5ؖz=����/��~~�9	h�d�#�C�+,	9l82,%�Q��=��=���s	?P\�Gݻ�d� 7�_n~�ŭ����N��ӧ'E��I��[����������ڤ{ �oU�Z������yT)�E������E6 $��S�4PӽS��*��Ņ^Ùp\���kf܇k�7Hd����6k��ٓ��a�˖(g,;E�1��T�j^k*�s��[�]�C��56o�B��֡�,7SL7��۞	7	s$�s��	O�ޯg� �j�����X�G�� 1T�a|9�k�!�H�6cq�^�́�w/��>�Y�8`U-�S���@�2d"V[��|����2Y��訐��ޥ��a|��2�H����ĮA���rw��,�r+˫����F�A׆�,�A��9�8'����{���@��9+tB���s���͏!cX�bEޢ�f�a�f�����,B��d��m���8=���Ja����D���Ӳ������7��jhض���ǩ�օI�[�Ø@f���,>\�t��K{��G�;�Dih!�����t~�����'I|4�^Ǫ`_Q�ľ��y�&�Y�[�z���HZn��(d��qj.�h&:[˴t!�dC��(��y���tJM�@�� [t"Gi��]%�Y�-���c���뷘��?�Y���I6K O�A'o� M��0/}�u�(��G/o:�!3��v3h�7����%�?,�}.N-q�j��m�8|=��%oP8�C_z�؆BI*]Z$8���Pg�������nfF���ϺwG�v�&�-YܲY�42l��8?k
6=�)�@�	��|֞�'D�]�����O $�Mj���H���)2�37�z�i)-���Բ��d�34���{��Z�l�̲�ĸ��;Ks�nߔ �����S�V��E3�❭h���@Myx�0�Ƣ� 6����V,�C��N+�X��&��{�fz��S^��B'��9�N���#��jbV�m�gk��b��N����@�(�+��]N����~Y�T�G�����\���;v,��WI�ٓV�k�7s{X��m��z��Ds#�����G��*Y�!|[ՒKCY�5�/��#vf���6�	��45�Jؼ0�p�-�� �iA�)xbIo�Gޓ2v	1.��Y�ހ=S��<���-��}�2����SqP�<��ȼ�j��q�_1�%�r]ì�2� �����Q�v2�;��K�cf��C�\W��w(��U���O�-��7�� 3z~��޶nd�=�#gk43nW����ޝ��*�P�n�d*���������J�UV =LǓf9���'��j9Hd�ƗwJ2H�:���`�����jDp�/�@��9y��x�^���b+q����g����]'��fZ
�o��o�V�A��z���DƫZ�M&^�"�XS�����[�� e�y&/�@6: �b������Y�9<б9Tj�D������Hv���sȪ����^�Q��
��]9��n���k��cpҽ��-�輶va�����`w`̾���A��j\�3��lְ��3r�(��1!3$�f+���5���>xEPg���v��Nu��,�#޸�]��Y��4@T��$�n�xA!�-�fD۫j�`�
%�<�N?�o�����v�DP��eMv)j����e׸<��� <_y���ŀ2�f;`�6��m]I�_,��0:	��t�k�'s;2�֣~�25r=�7:����e*�;C�V6��R�*�.�~Ew4���Sa.2!�q�:�a�i�͓��4�I�$+� ��v��%�1\�r�(���f@�(N#�,}�}�W�`K�
�HK<���w�+I��m�<��rP�5���W8�7�zGI.־��̡sy"K6���7�`b�>�eJCBL�RAXn�����}Jʂ��J,C�.Ǽ�!���Oҭ<��
8)vA'`�,e_8=���%�]-ú�
9;X8H���+{���_S�'�R�-*�cp���(����N-�=��W�$UU��B�N0��_g� ��`�D�j�Qk�$�\��ʹ��=$کJ�_X�C��w��{4L�h��j��j�Q\>�1�K��m��Ǐ�`(]=\8��Q%�lĸ���"�J⹄T]Է!X��;��r��R�K8��D�=i^,���!��,�#��P��X�A�C ������!������ib{I�/T������f9�� N���&��ҡk	ϽָXcT�|{�wD�>9�d?Q�fC"
{��.&���UG�=�#7���dʎry���\Tl��ȫ6����5��`VR����0RE�Γ)�ꙧ�s�ײ������J�J�5��������b�(�A���d���,1�/���PB�n��U�|�2g
���������,>�*I:~����ٵ5Z�e���3x���ƴ"�lj��w�`BPg"$+�O�I�GB�f�<���F%b��U���u�AFg��T�C3u��+�FqWR&@	)s�.����j���g���!�,̊ n���@���#�v�؆q��-�"C�E)�XŮ2�Ho�|6Pm��'�7�s�P���͒��EO�8���s
YF�T�'�S2�/#{NE��|�+������\��5#¿��K؀6�r�.U���6�*����v�0�)��������Q~���E��#-ɝ7F@�&CsLB=�Ŋv�W�b�z*�i/�b�x6 S`�R|�׻��G|�-S��C�DC�9�bL��+�'�2�� �}��^��<��*��g���Jqa��u[�����(��%C�?8�Q���� !'e��S�����/���(lz�=��K�����4��v����0cϊ��C�\s�8Z�?ֲ���^c#�!�aƼ��~ȥ�S�E�+�,�<nj2/N�3,#�k�^��٠�++�Bg�C&�a���ySN�$�L�}��@C�^~�%,	WMFk�m
�h�
p�K\�ʵ��o���������ZI�(c�vN�+ށ��F���,߰O<�g�����n�H��:��զ�����lso�F�1�*�ނ_�H�5MH��:��O���v�a3,��V�������#[^V�u�v���W���er��E7��j�|}��C3���"#"<\�����s��o��<c}.���1*���;b� �����=�uU�UE( o���t�!�N3�<���_���]XT��C
��}�h��{�X[ՄM?Z衒*�2��L�
���y?r��]�;�9qKmU��$�sqqI�(w�=�}P=��Z��H�jq��O����*��.�B7��p�`����3��.�d��i&��x�s�f4C�I�`����m#���uj�����a�ǚ�>���<ҷ�H�����mM_�'�C�~��1�Τ�O�ŀM��gD�Rd#rr�	Y�-�S�A4��܆i�rEr}��ɼ�h*Wj���'�yn���:���[x�;8s8\0�xDH\�d��j��r��%-�/�Ȱ{��1�t�S��2��c��a8u�].��á}��Tjo����֓�R��~qk+�(�H�{NEk�٢���?�6[��G�|��:3���A/��]�.*r�I٧w����RkhD�9�ժ
1'�9g.3����e�t��?��������b8��iqH �/ն�P�<b�܆�	��Z�Ɇ��=�P1��@G��6�
a3���-�� p��+a^��oxٮ��,Ƣ@i�u[g=��[#ʉ��&��f9�:P��r ����;1�I{�h�$��w�k3
Z��9���i=b�_�o2Մ�#�X�ǚM3�3�2ڡ�{��\�t�Q�K��k��*w5Í���aQ�q�Tt5��E�U�c��ѕW�1P�\]�a9Ǔ�!TjG���y���E6���[�+kZB�-O}	�skΥ6n�H4��l|)z*�E�R�`�s~6�l8���0#� j���n�p/�����`_e2:_]���+���0�qM�;��urK��\�ϧ6�:+��}c��o_�m����SvD0�_KD�Z��) W���X�]��њЀ�Ķ�	�x.���_��i�_���Z�x�`x�+��o�&�bه�_ �=��k�1�������y�B�U��FC����#w�-�d
"�����ͪ�'X����K���UF���d7g%;���Ac@�hL���X��H��
���!��85��!�~`�9h+!���CFO��L:���o���r�΂��l U���������{�=�j'��uo8@�=3e�g�k��0�x��Hڰ���w��u!��%Nx�W�Hj�����D�1�����_�����x�f����q@����!ll��i��h���,s�e��Z�9��Ƙ�a�T���^�B`�ih ��G���U��H��3u&T���%����x�oe�Xnkb�#�������nln�_�s�|Q��S�?S��t�yU�i"���T'%��G�wD����fީ�3��"ͽ��os���]��lX����x��_����]SI�^XX�=�iuOG�U�!9�үA<ꋀ���?�C�E�N�����N�<�OYqI,��@J+�(?0�S��7"�~�y7i�`h��SI���26l^����oB�	�,�vo��,t��/��e�`����&t�{�� f�4b=�0ֶ.����"p�*��_�Dh�W�qN|T������ˬ�9-!���h4|�[���!I=F����"2Uz�0���+��YԬ�$za�~U�Fkado.c�8p�T(Ʈ$��%�tjw�����t �n~��_��������&V�E�(�x]'��אoY�M-����F5ƭnbp�e�:��|��gF�EHuU�O�=����0F��o��%�g#nI���,T?ۣ�[[BNW"�E��{ߩ�C�D�j`{|!�O��!K�F��$~�Pi��ЬK���`4��)�k��J>�YX��[�|��˻h0���sb�-d5��6�9��S0ل},��`5�T�m�9O 1�{��4g�Y!T�!��9D����*o2C�վF9�g��lKV�paER�d$��Wm�| z/���jT�1c���#d������g[���.~�������Bl��"d�T�<�,�P Ma=�X��F��X��/ꇰ���Ín����1������jf�ZՎ5x��c���aX�Aث�O����/�j���>
>j���p8��{��K[%�`n�=�� i��#���)Lm��K)����\�f ��Qm��za"A�W]ޖ�|�}���FcN���ceP��"S;i���?P��v��5���)���%��#�  �E��4%,I"�:���u�)�[ța#��`��2���D;J��&��s.3�� ����Q�����ݼ��j�\+�@y����`ᄆ�[#7	m�c�i� �2gd�K�o슄,�ą����x.L��ے�#��9
]s
�S�9����z�35I��XW���ާx�}W�C(�chX/#Nә�i _فsf ן~kw��\�Z2VG[тUѲs{x^��[ًПq�[ыܡk��7b�~�Z*�c&ԙ%ͳ䁛/3�l�s��i�[���`�}�#����{���P�H�r[?|Vչ�M
AB����������	���c3��W�I�t�u[ab��4G�͙E��3���լ����� ��� ��Y�''�F*2���,L##U�`r��ޖظT��jT��Ee�r1�ӌ��Yl{\8�F+�Z��Ƅߕ
�t���Pt'`��!��S���`^g�>�~��0P�&���_�q��ֹ�P�+�>\�a�h���SA�]/����;��W Ⱦ�F�нǡ�����k!-1#��& �f
qlL$�`���0r�^�@%L�i��	�{b�y�`� h�I���:��	�}=�
fݯ����=��"f�c�V��"	��+nV����X%��񟸮�a�F.�	��_, �͔9�cL�������4�H<������w��Fs��V��T��oM���~w��p�� ��ŀX����`�ƻLkv��Δ?k�?���"�>�Ŏ�	'C��W��/x�B�\�%g�����
��׉��:-�$(�Xy��^�3�#I�!~��ׅ���dܖ���I�	5+1o���k�U�����̈́�9���b�d +�����ߚ�X�6p�� v/'H�+�!�]	;ˊ���C��gR�*_���h��|� Ɵz��=9�~�y#j�Ə�A�!Ӕ�lDEw�{��6��)h�\+�Q��l͕�a�^KJ��釂�Y��xf�=�53͕J1Ka!���P�]G�R{e�l#�N�����0lFs0R\=;��8ٸFh���w7��=:���`A1 Z�ermWZʓ��?�x����&�m��@�)_L�I�-�,3@pHYt9��T�8b��{�a�v�D�W2p.)U�R�נqKag�0���~�SĖ��'�y�xL{�I��6��;X��"�z�n�9f�a>�3c���vϋ��F���mR���`s0����y�j��(���f�6lft{�C9i��1Ia�BT8��]'�� �̼���ɧ��ȓk�v<�s�k�������J���h'sٞ��<g���>��<>�ɲe��8f/C��H��*k����wo�	�o;�/�S�$��eZ���L	���o�,ʳ�tR�g�\*E�J;OG���@OF��0����`2�[f-u��0�I�*)�/���y9A 	zp-���̉9i����B����V�ô���"�p��_�O�/	��F��\�W�3�x�y �?è�1����u|����������Nn3��N���s��aPx��y8�w�:�K�^����B�#fo���Ѱ�A}��@��xϿ6 ~L��Eڪ��{���R\3�cW����	h{�J�}#�İX�V
Չ�oBgg��(	���yaM��kh;��J@t�y:�p�hhĽ8F�� "�$�N��8�޴<��Szrsw.0c\*�#�$KD"^b�������D����.3�ǟ�ntc���3������B
u��/5"���.9� d��N&�=P�p�y%&�z<큄�xz�s���Y��8��4�|�.-��&&��3��)��v�m*C�P���L�E	����q�������!X�R&x�f\CL��>���y`���$9����`۶����M�{�Fkh��-O��븚��.ّ���
��K��-O�M��?;��E��:'��1���/8��m4t��"�Wh�����$��N{z�0����G��`��i��z&�0R*�֮KO:��)�d��I�Pz贞�6�h�Z�!Y �,v)Ns��9v�F-�z�ַ�w:i%"�e�#	�5Jwu����,B���R�-e� ��Ԥ�2{�I_ͪ_(ٞJW �hd�GG�T�Y�E�~����P����e�Z��p_�G!B�W�a	Ac���3X1y�q��{Ч2��=�9Y6Of���[���Zq�X	�bZX�_�S�!��=2�²x;�^���jj�Y�ۜ�)v�Ɋ��40:e`	���ĝe�<���1��X��mR���g�)�(ʔ�����s�nî�;�6,�`��1Y|�Nr�Z���k��U"|5q�8K�����At
7�Cc\:����lh޽�ф�Sd�3L7n���y��uJ�뫨��"��J�����G]��h �M���C���SÏ�X7�Ȑ�;�n*UT���ةc�h�/�k�Y���(H֒�EP$E��^@x ������rl��.��_�[�S��ñ��7��q�[�04(�b�2�kw�CIC�#�썫҉���[O�x��ޣ�'L��|RW�W��t}�@
{��Jg�>����6Ѽ ��7�]g�iLU�7���D{M��h(�`��=�O#}FK5}m��	��e0�2{�)�*R��N��=�m�Л�H]|(~HI4��#�[��]6�&|�^40�v��#�}���a6����4o�h�t�$��cu�s�0���7=O'�JC3��O�n[���n��M?����x�;p� �4�pm�y�r���Ѹ7J��ȁ-�	�m�͉���z�b_wiI��I��y�~0�o��Ys=#u1sJ���}žJ��8�$�K#F��=0�x(l��.�<���X#���"���N�8��p �g�rJ�e�F����:�y?GyQ����$�2|_�Tԟ00�i{>��g�_|W�Vv-�H�6-]���E�
`6��@�������g 'k���^�n�lI��Rhinq����Y�����F���b�X����2�S*w��@���j��6,Cz��K���u��.\���L%�MTL7D\����O���b�MG�|=t�@�H?����p,#��U�T�D!g=+tiA�_!���,��4���pL��6�*zɐ;��d�e᷈��Z��*VۛI�������c�G�׫m{b�����y�R���)��4q>����`n�y�N�&��C�E���5�>�Q;������w��_��z6%˞z0?�z ~�s�8��ɿ�d���hN��:2/�H;}��a�Q8W�����nJu�>	�S��T���p���LA��=�����-�-k"����:&��F�|]�D�Ȋ1����zRd����Db��ׅ�����
�*D��"�Y����h^�͘�_�����L}5VM��]f��TW�����F�]:ڿ�:�=`ze:�[Z]����$�l���,��^�����Ob���K��d�@N�-��/�M��'&P�\)�s P	��M�x$��U\��:��<Q�^�ܮ<U=��N0?XE��Zw�2��aU��>������Ґh�CS�����{<�L/1�ɍE�Kr'!�7�G8��,�B���Z���(�S�л������C�P�hO�U��"!���xkȝ46�&�ƩН<:��$"�{d�������$%1�$��`+�&C�䥧'ޥ<>�E��`GLt!:��S�Ue�U��Ӭv���?��y�.qX<\��̶lF�#ߎdN��w�,�"^���s��'�ngeb���������U/�*��+�i� fP����2	i����?#%nIbRf�3s����cw�&=���!�G�T�W��!�C��yhZ�yw��\�f��٣�7��o�N����A��ɸ �
O@la�C{���,7��-�,��ǰIk�;�J4i��;X5AMԋcZuw��
ua΃MX�r�,g��1w��xji���n����=K����4`�v�U�
��o��D6r�J��Wa��Z�p"�or>���%!�,���^����$4?);݂V��x0��k0ɰI��w4m�ǌ5�;B�fA�f�P�\GqU%���i�r�.�H/���τ�����iǏ������;Z"���WX��'��r� �zg�E�\�^j�ͼ���.��x�2��&"�����O&�W�R���7����f�5�d��Q������߂�"NJ�P�2ʺ��>ac�4(�G���hVQA��h��r��s�f��-x<.���<�g��gS:�J��+5
9osⶸ��!�L�&�RD2X����ǩ{�$�cϘ�9Э6F<4{���Y�x���/(}*��l3i��Z�3cx>'�z�"�l��r7`��~ f�ժ	E	6��.��Q�#b�z�2�j�_"C[��\���=B����x���r�|�|R]\)mw�Ta/�~Ji�@zE�\c�������r��:;o�Ʀ UrЩ]8��h�v-ɵ��mt�# h��t�o�L�-V^z��H�>9Y�Hg��^�?qd%� ��ר�65��	Nh�ٕ�3l�|i��D��K{Q�w�Y��CU�{�-f^��^����F�,n*ƈ+��&��mG�`�+@��h�y�,VF�₋`t����'�6�i�����@B/��~�61M� �1䟠݂�e�O`eV)��&�35�4����o�-��[�Sj���R���S�PQ��|���,��2,I~u�q-�W �1~�o^�`�Z�ŝ����+IHLO����)��, FA�~���~��]Q�pE����{a�?l��(��d ��%�f��s�e׺�Rwf�+p��̶�3G^~m��<2��`O��$8)}�L_������j��pb�H�J�ǩ��PO�/�d�HUw̑�D��s������&�}5V�@|aU�	�ے�J_� ��4G�NFQ��>�%���z�����]��1�ي�՝�Mͤa�D��(�*��_ɟ#�F�Σ��D��s^����T�t�b����6n�0ᇰ��U�	�Ì	g�f�����QB��ux�|[�w,oD�B�3�xY������_=�Sx��P���W�����Q`w3#�Zo�9�8�"X�����q���Gl�m7<�e����/N�4�%�+(��e�P��B�+?�����m*�S��|%�tZ=>ёq��u�u�@���0������S���K{';�3����jCѕ�����y�Y����w�������{��U���J��B�hk׵�ѐ��%��/�h5����t�?Q��Vm����Y����4P�n1�R��ML�8����gF�i5[���9�\���/��.���O�M�� �o���uos���/j�,n�F���i�=��5�*ǐw#��#�-�2���e;��2�͵�\PM�"?�0*&<��LsϹ���H����h�}��;�C[������m$�ُK��<B��"��QRHg^���\&J� #MS���>]�+cm�l�+=OZúbUk�8Ɍ,H����%%�xb:�~�
a3k��L�~[��E	��_>˺���f筢�9�,5(��v[�ܕ?�f
�
���(CC�0ou���7#uV�̥���7gNl�b�:������n�s����E��*�q�G^X����?[P�7�vVVy�1�C���=U=6x'�.�a}u�t��<���A�b�3P֐���%��Ϸ�'�]��D���JDԔ��--�oħƄ w��1V�aNE{q�����F��e\�j	(���M�`�[�u����+ioE�Se{�@y4�Y�ۣ�3��.�f�<y���إ���z�l�$+P�Y��Y� �*IGp,+�|���~�X�����>EV,��}�U��=�kR����:�YҼ�z!�V�^�� �0�~�����!#�ؐ��P+�}����I~mk��
i�3.k�u�E��ӏ�52@�%����1�y�B:O�����xy��_&@\d	K��RXR�UWS�~G��[��(#J�rB��h���pT�:˓�������t~�,n=1-��'�T�Y/Ӌ
�]�����Wf����z|r�1�*p n���XHP�xx�$	Fu�Du�>?�.�ȥ�4 ��&�K|��l���O�g�.YDor����0��<��ͼA8�M�X��[�=�C��.��Z��z�A��kG��}�a��V樸�9"�W�N���_��k���X�+= �e(L��'��/�>��a�/�n̍�%=��MکU�h�.��v)���'���	���?�7\p�2	v�5f������;�u,ˌ�~+���»w�:��Ҧ/��;b���K
���ͬ.�-���b�#�.�ڒ���	x0�6��E��Mk]�)v���dv��(����$����֎�x%
���s�����N�{�kaY�n*��ǀ�T}Aq�(�����`0�5�ѭ�R��;�D�j�\2B��������6�ASM<���@���soibS{���'�;��=���P��v��xx�-t��?�����"m=�[���~1변/?����X�i�P�H�C;�d+E���h��8=�9���^�����<�"m�M��;+�|�cI�E}Mc�!H��)�G3��G�>V�mR4s���T�&3N���<SwH����/��~��^swiR�9S���ܾ�eE����(���f��(���(j߱CUM�䭒;���6Cl��?��㵷ũ�)fJ[d�6X�i(��r֟t��T��������7��\���]����C����P���)����
d'f�Z=��p[�Q5�w�̈́Z{m�x���Pb��7����Ի����}��3)F��qH,`VŠQR������皭�RQ����e���i��{��	�h�S��F��&mĥ,^�K#K��:�1�F�[�:��WE�8 a�
g����-�BpLms�9�3����o�/.�ەǍ	RW�gRwM���-�,��a�|�Ց��s_�suC�3�B�i�u�˂�o���H��f<�����������4����	�E+Y~�z�_C���UQ�M䕴����aK_�����{G��x�bt�!�8|O�]�^�!
�������}��ۜ�f�C�01ǪE�?�*����,�Vz�e�Z\ϕ:�C���ӹ>��!S���X�6�?ѷ{��R�=t��*H�p?(GQP|xӭ3	]�`.]m-���.��~ܿ��C���Gf^�rd�|3�'�擺]��(�4.R�i���G0�f�8��'�g�@���A�.�q��-'-�g)"���0�"ҵk��}ҹ)9}��Ζ�<Hus�Ȼ�e��,h?2�������	�Fb�wa�t	�Rdų�J3&�9]�}��e�vԠ����c-a�7�f�^��3�Ϫ=XE�>�{���l𔹿6�@�D���%�c�4JExA>1�l �����k|���~���R�޸;]�2��*Gnb ���*��cI;-q�K��`��ޗ[��h���9��=j�0"*�E7 ɫ8@�T���H��g�p�*�P�r06��������ऽ?w�����+4&H&�a��ޡ���h���>�k�^!?��JJ�K�������A#��8/�ʷSn#��4�z��R[үκ���ŕm����r�����[�<�B�D@��^�t�{��^�e��K�F�Qw���oU ���Ծ:A|���Z���\���P����P�������ߊ��Ԯ?��H����FJ�!��C���A�\J^R�"r���]��]�}~��`~$�Pz�T�[ʘBY��'F'v�����6����O�!�\f�����Q�Rս��댴��ю��D�)E{�6ļ$Qy���K�78uo- ����P�� ���4�!N���&�#KOS�T/�t@X>�ߔ���L�N��	��+T�r�H��P"����ep2�CP��7U��y$P"�Fa�R
���e=�8�����"3��o&�K�WIHe]*4-Ď��'��\)=ϓu�+�p�Ô8y�߈즰��mV@{hْ~=$��p� �b�-A��N'i����%�������b����1�E��q`?@ܩ�k�S)z>�i!y�v���5�#�B��k'��3돌�x�x?��ݵG��찌��˔|�!��~b�ψ4���'���*�^����Mj�����*h!�HL�Bl���ɗ����ˌ99�T,��\&�3�R��Y�X�<t� _ռ�º�hS7�}��X���NqX�f�Щ���J�(��V�d42
7��2���2&o֖!v�jl�sF+�]�/��u��uۯ#S���*J�'��P���dL4=É۬F��P�wK�����F�v��[�<�Ae����s2t�M�Dpڜ��[)I]ŝ�zr�~�����5�F5&�a]�歏O0Э�@�q�-��D5, �I�3n����{~�oc_zN�%�X�6( &�U]��Ug4���C]'D�ц,����m�
��ӭ�X����d�W_0�]v;��I������qpЗM��uY����>��"wچ�="b�%-B���'+
��q�J^k!�-W��[/�8�"d`l2��)�]�R#����yf9���k-k�C�믿`��<�� Cs����ɣr/�>c�ܼU���C���38�x�s���'�({��p�{����!�ց�wv1Ƣi�8�S���r���㴶GɁ����'���'ĎP�ֆ�8�(��@>=��LiA~]TF|K �s��ĥ�R����"�.�Y�].(g���Ib5��9�K2`���m2Kb�g�C�?(hp�l�dn������p�[�P����2�h�Ɇ�����z���)T�)9.��g����J\������};����<Lx�r�"�[�lQؙ����Y�McrG#h�g���{�Im��7�ߪ�ޟ��=���N�(+*|��׏���>�Ķpd��ʷ��O�n��"u0�� �!N��4)Z1ݘ��s]�ppxS����9��]�,:k���"F���Ͱ�KD�7MS��n9����0aؽ�6�$V���$����,���_��Ó뼅��I�?���\�-��#�����RLPv!�����gx�A���6�qb��L��rB��	��KF�$���yM�7���p~�j!��A�6�����^;/�v�mq�Ai�>l�U��i��,��V�[�n��(�d�^��]��x�0�%��d(ӌϗ0h���i;���A� ����+~a9�Гh�I�!*�<�h���h����̈7j�n�2r��ٓ�dM8���[��k~e��� G�	���>�k��p�� h��E��l&0���]�s:B��\S�f�����2ʦ �;� ��=�'�����p$Tk��*D�B�ť��/���8�=�K�u[M��%�q�m'<��c���؁�@�_��M�Ώ1~C	�1F�_ZTq��p:��C�gЉt��~������#%D���]�ć���P}i?&Q\ggȫ�"
�ԓEF�!�	�̷�?��Tt��E��e->�'�y�(
�B�L��|��Ŵ�Ş��,�Mij�fI������j#6�_ED1~��p(rU���<��t0�9?�a]��)@͔Un���a\ĺ�z2����~"샘sf���S4��[I�J);���ři�u����j1౩=�,S⩏S��۴+�Y�ib�r_����p��#�M�E͝��~��JLo]��C�%z��V��Si>�w��vij�s�,��o*Kun��k��i��������y��6���~� =��0o%
%��Ʈ]������TȈ�E���!�T����4ժ__��%M8�Z3���ۀE���ӶE��^�!MaʐKVR-�w
��z�E��� ���|׽u���#��V��ή�3���}���/L�b��ȏ|�-��Q�H�۫�~�$&�\�:_��S6
���|$��NM��]��l8βK�GA�t. u��9yل�w���eך��!w�Y.�+*O��&����N�k�	Q�y��C�H�|1H6�a~k��H�36��W/*�^W��mKu��4�`'W��o(t��X*���d��e��L7\� J����}3>c������� ��ҜJPe%��٦q3�C��ҋ�Tj�$�n�q�%�G.�L�3u��A�.�)d�����Ȩ��(�p�XkEIM8Y�a!]�<U�Y*���W>��tJP} rǧ	� 9Q��l/�iƖ���Hss��z���.i@�z)�tϸB�M��Eɸ���/��7f�>Ҹ�L��li���(�"����I:��~��A5�����өoN�@Ƃ]��3�m��FO�ӎ��eT`������Xj"���C�m	u�J�J��Zw��r*�ރ����)�b.�	������P����cw�\�i��	�8=�deWt}ڦu	���>/z��NNܲ,�+������'�O�ph�O�-�����ݯ�!��}��tf�\Fn��M���tTF��������,Z��V�F�����i�*���+��N����+G.l��0��;��`���ɣ�w�������q����@� F�V��GM_e���eV�����+AV9�GyG?�!�A����P����|���X�c��_�ah��;�ߩ���>10�|;1�b2tw�dr��YC��4�~cbѹvY���&ЋA�:jSX���h�!��-�P�V�]����`*��\�X+�Sb�,Ǣ�4d[Ц�l�TxQ��)߼�i>I�c��z�l��&�����{��$�{me�AX0:iFLT�D�m����),��Q���}�f�ٷ���Jf	������U>U�������3�ۭ^)�g_;6jt~����-�<q�h��M}�j��沝?�8��w���m���::u��9m�����K˞)k�Y@�?��t���,�|�L��vDE1�b�:��1G����	�!S�6]�+|��@�{}�X�D��Wx�����U���i����Ժ�y�9^xAo��,]����-�څٴ\�C�B�l+@OCcqQ��iRAJOd���&]�����kJX@�gU��u[����
��;Hl�qF3���az�q٦z�6G��p��-\nY,}�RW�)��4�cX�[�2��q�la��X@L�\L�n9I�N���TW̪���
�~b�9����)I��Ƙٖ����d�ꌣ8=Ӷ�<�����J�t)mM�] ��x8e��q�D_�+I�`-���t_�*j[BؖH5{�m����s��.�Ո���#h��5�
X`�2ț!g��]� ���\.���!�&�ُ��+�z@���C,R���H	���
.��Șzj�����ρ���D�#j��G�~P�Ɩ���o<e������D��d�o��y��iӈP�.d5l���֡�~�C��7?e%��m��wx!C�R+7$���٠�L7���`���o�L�emqGRhI#��Z~�"��FnnX��o�1���߹��s����/���7�'�6�j��?X�����l�i|kt�˘E�⌗��mi!p��4�ѐ
�5? )#0��)F?0���n8��n���$(��\}��S�e���ӽ,Q�9F�*.B��(.�t^�F�0 X��U2�����;᏶ݣ���U:��`	q�0bu�>%JO&�l��F�	-]����U?#�N�]�*бS����xľׄ*�d�]d4�<���`ݵG?$���УкC�L�Leu���)����#'�r@d�U��;�M�^�8�_  ������I�&����6k��-�/bi��.7"�試�h㛰���ވ�c�h�Y����;}�Q�`�։��̈4�/�@Rvo'�ڶN��nb_�:�TCMⲎ�I��=�����.�U$`<g���*���i�֨N�`˧M"<���%�FSW�)�[���X�/2��J���?OW����P�;�"��7�?�@���݄Nx�|��%�	����%AC�����q����޼w&����w��FB*ϵt��|S�-^�U_��jI��ȗQ�ģ(�0�G�d8jU���)��F����Ƥ��p!}x�V��H�4)��� ��՚Q $�yϨq`��.))�~�X'��t;���Sy�vS��֤֞�Y�L�NYTa�QJVBj��}��QC{�z<��2�iK��f���o�u��m��+���y
��<E�_������(L�qM��@�#��Ύ����-vvE�\����S�
�>�$'s�cL}��G�Ȼy���v�䊫��Y@�"���y���Ӭ㜤�EƁ�!��(?����b9��;��c�a�ä�bh�NB� {`x�tQ�i��&��7�{�Ne"����)Z:��.9�9IJJM�D=7;É�1�� �'r�KRu;YS��EsG��G{��ֲ����c2l>�m($����w]��(��Y����eT�c,�+ �N%�0�p�Y�M_�v�����	��(�Σ�߮��4c����'���
�(9xD:��OU�Kz�AvAWU-�����dͯ�0B���{�Pa�Vg|�K����W�/%bGw/�3m�p�?�f�~,�l�����������׭%�w��������R�����]Ÿ��˛(��cX/�g0W���}_f���͒������wQ�~������Vae��N,@!������H�*H׎�x/���
�\��|b��0�D�Z|:f3Y��q�C�4�f.���o�)��#ԉG��{�/��� �Y�>�U�
�#Ʈ�WL��[����Ցȥ�8�`ݳ�k�]Bx���Hm���~�S�m&M��1�{�0��a�ȅm�c�v��{�۶��ח�7�p�=�A!\����<b�e��b���S
��Ap=S�A�*�b��m�Zt�0De���z��^w�����>�G���J/]=��O �0�#�w�(�-�9��� p=�Q���5�>V+�󺨥�^��ę�{jGf�X���1����"d\��?�M|�N���G�}e�5�����b	���OLEFe�&!Pκg;B�lH�^�8�K!�#)����*JON��6<)�&{��a��e�f��ȭ���Ur��	Af�\M)��n@u����ȗ���x�-z_�����xƞ�;z�=��`���g9cf�x�-��� S��\��H&��۔�a+�=jv��A�1�ֻ��+ʐ�XQO��J��a�����P��g���6-L���D��<�הS�Yn�?�!.
��(�8��X��e�n�x
������o�>�G�L��gZ��A���xF�����[)�
V
��m�o�o�\@�3�u:E�?�f/��7��3�E0��f/�D���l�Y7~�Z�G�̒ �
ș�,��{v�g���g�bIBБ&7n��j5[TP�c�tD��P֚��#mE�ب����U��s�7�=�͢��n�s�žiY&KL*�q��Wq��]}��!�*�^^���R��qp2>�
N{�<�QV��W[j��&���z{�#��qQ��,SHQ�8c�LG(j`��pr��T1 �b�b'8ù��n��\�����6�n�5K�$����A����5�Ζ�,��QF}��� ���}dE"T��"�-N��ݦ�'+BP���H���d,���]%d0�=^��c�����l���Z(�a�/��i���Q�H�)q�C���Ɉ���@��ۏ�Յ��WΊ'�6�e�m���ñ����8i+>'�W{w��M���y��d���2֐��;]� UFl�ZM,ÈN� 	Y1�6+5@'=��(�<.�����o���i����ō53^b�K�m+��C�D܌��10���7����	6_��]������=s"E@�~���D������o��e;^%�Њy�	�R�WՇ#`�N�h[yL��%WK�B�I���0
�~�C����f�`k��]�Ƙ(�Q�9Ǣ��u�\X� H��ɲ+�O_x ��%�s3sm~�Cc�G�)�݉�e��h?%���k�@����|�)M ���G=z���_|��x����Z5��5�6��ݏD��=e���W�>N`�	��!����)��Iv\�v[ ST�i
=�D��P�:��{��qp�孔���E���?��h�tIv��Y���o8�īs�5sy�!��7������az�Ԭ+7�����3��3I(�`���G���8�Q�}j�h4f��J�|�]^�?K�sV����s�*�M��	�lxk�3z��p����lp���껰�N��2��-�:�s�[&��\9�����߮�9��H=�t��7�)��m1W�suDoZ�)�RǨoπ�W��L.�K�LU88��-v�b��SÙ-�Kϙ��B\!���v��hEբ���I�-]��U�͢<
�Y�zIrOu�v�s�L��gJ�CG��8Bm���I%��nK�m��dp��3� �e(�U��z7��躬��Z�F,��}�@�kv��v! �6��4|i��z	�-�.=�ɷ��8��6�9l�ҕ�mX?"�ql��5)|�"�k0r� @���H�%�A䤸�a9����=���׻	�1K����Vy��y>'p����`Ol��NCľ+Z�1-����h�U٨���D�F��(��F�@PY�V1V	}�M1wV�e��O�M2��g�%g �.YRǕa��#�V�o�D�$��u�V���-w)1��
I���m쭤z+�u~lG�"�����vǐ*6�K�h�J�]�{a\�^��79��5	F����#�J�~���7��ΛL���۱ñ\���H����c̠��|���QD�p6q�Ϊ��\��8�*�d��Ort�:r��D��|���5m�#���M�`�"��b�c$��H!�xA?_5pf��E�ߩ���E�YJ` >�<���D�����b��I�~��84�.�s�@oU�~;U/a�ߛ��/zN����azvL��hX	q��Oj*W��ub<*Y1�����������XaEGP��ɋ�[�j�H�b��4F����k�X�?j��
�С��2��xP�G^s5U3�2Z�;��Z�H8n�NY���د�3^ �/��R������bQI1�Tle�OK��a��%��{��6��Yy���1���1��
�s��j��6�nc�en���P(�J�m�~,�M�/�C���/P����
�/��O������~���6d{�1q~̺�+|�5d̯T��~���{�}��0���%��I����Uuͽo�u&�w�@^Q�Q�Kf��G�p��'3���"��+2�1׈���m&K���P~<�N)I!&��n|C3��/��;wp-���27xn.]�>�������˃�/�of�LI&�׭o�4�d�`�ġG�����Y���i��\'���D+��g��E�NcL���৭S|䥛AyL(,-�t�M[�@ t!߳j�-l��A��M���Ҹy�O���lH���^ܠ	b�,�#̔:rg�������N�04� ϧXX�-1\��"�~c0�&��k�5�<ʁ�O(9P�c�6�f]�-"w�����x�{Iu��A�x��?��^Ž/�i-ڹ�BA�"�i%�N�3ύ�X[Ѯ�]�7$�޸Fk��ٲ�`Q%���9����-Ï��V����4B�d�m���k/�K?���c"���'j	����{���z�
NƘ_Gk�Ow���rx�����u��KE�����d�L�P��m�5��]�]z@�kl�lIu���D��B� `�y�J$5��W���ޖ�}��^��k�y���Q��m��k'u�#uA�z˩����@�`�A3i������Ys�j���a�oz�9�vZ����{n?�[d
����!���Οk�Q�Q.�S��)�L���+[B��::���%<Wh���^~���Q̌~4xg�XC��S�{^�}���r��)nT�u�Q�^�yZ�᷅�SG�9���r\�N�5ձ�x��k&dp'�Lk.[�D�F%;eݐ��n"�����C.�*�I�Y�0�:���n�H�ߴ�&�>&49@!Q|�m��s��bC�tOh�Ԑ�$L^��)
��*;HV���.te	 n�����f�c�n�� �=�8 b�8T�<��#{���Fv��"�j��䪻y����y�w���� ���1����	lU�l� �u�ad��8�Mf��h8�`��-0����ņ3��k�8�U���u�)��1�ĭ�_���_y����Xz� 9
�Hk�r����3��,V�*�-��7�Ή���	[)C�p��%�Qy5�����]9vߪ:��q����Æ�����'`������j�Ԙ�ǷW_�� ��z����Y�|���gY(�9)����@��w]]�Hߋ��Rf���X^�Y�-����7$��5�a`a܁��U.z�n5KB�/,Z��r/�'G����Xm�),� ��Y����TV֒x5j8f͝����fǣ���_'�t!kΦu� 
90����ʫ;�/ΧQ�G���X>�?b�բG��8a��[7���~v�/�=Qӑ>	1�G6<�Ꮉ�1	����C��)}�n�Pv����;&۽�0�E9'�R�bB�pO�w<E�R �����͂!�):oL�ô�.Ʈ���Z����xs$��=BI���,#����\?�yНR�bH�ƩC:�s�e�#I�4Q~��\ ����L������։w
ȥsIuR���/Ŏ*����R�J\زSI��pE��l��@�K!��W��4�!�@/�gf돎}q��@��E>����D
�h�X<Q�-A�Y�v��������<:VS�-n��Г�G������q�bű�(~c*��av�R�Si��Y�ż_�p�f�j�(�.l���]���gȎ=�Q ���;�A�#�?���%�{��j�S�(��IO� �Н�蘒�,����N�}�zL +�����u�ܛF=L|\^K��XC {��0{m�Vr��`�|���a����v��08mWg˾$[�<���Z`�����݂��Ҟ+� �u��E�| ��^߯�����݊��$;<o?���yj^O�]�_���*@�ޫ�)����g�?h7�B�./܁P�Ze���������NU��E�F7LH3�^
���k锖_��jہ�@��KE��J���]V�N���}��){�G0��V(䐎�rE�u�E���Ûض�{��*y��$��"��×U@��!���Vk@����������7���(��� ]ߧ��>��Vt�����^�Y�4�%&y�.�uG]���#�NT���=)B�,���w��,L�b�����&|�*���Ⅰ���'m�S
��~�/����E;V������kdun�..S �h�WSV��+���_�Emxk@���;W��0g�<�hw�9���s���ƚ2ѓ����E �ō���?m�4P�6��@ƞ\'�8,P܂_�h(�2�]P#M˽v�V.�+W�W!#F�C�����C$g:���T��J��h�>����>N���؆,����R1���/2��A��N�1,&��4��p����'kn�u}:�:llR@�=A��c!}+O��W�6اIyy���>V..��riR��o��CYi�d�v�NkĨ�����'�@��Cj�@�� X7=�:�q��M}�^����-���8���|�s�JVȺ�z��x�&D���MV�{�����Y�EA���D����J=�lS�Cf���x\��m0UE����ZnF�(+D�Qg���8�
s}G��]�ͼlG���mF�'�h��ըg󲮣�1�	y�jݜG��pDU���7d������AG~ֿņ�ۡG��#��f�|��~	h��<R+I��M���1%��
��4͋J8�xKׅK�O�/r��>�m�&*	�%��O��{�8�NLL�_�KAf�jui�"5��ܜ����O�g�4Q���7Ҽ�よ�b,�����.�z���<����ԧ*$w+���^
$���@�)݅<'a5^��Z��X��,�bK$��"�qi��(:%�{�4�#�E�#�]@�w�i����&*jE���^
|8�F 6TݛȘ�Β�f}A�

_�P
�Y0�dxi��:AT5�$�/���ܖ�&x��N���	�H�&7'�L�Z�/��%���r�!Ҹ�ioB�����%�H��g0y�����Ď�r�aF=��U�	u�(���5�t(8Tb����fw� %`+�%�bM cy9��a
>a¹��3Gޚt;��&l0����t�ZjC����v�Ƥf�4cz(j㜔�6����@=�r?�@��q����U�*��=_���+��]�<)8�L����9�p��hba�eؒ�q�5�v���b�����KhM���?�')	�$`���i�-�5��Fjp�=��n{jQ�Se,��x X�c���s���NU�K0�$Y0����j �஄�-�@�٤|�E6��C>^O3����h19�5A�]���gb�G=a����3������J�wTbW�m�aO|mZ��ꌢ~AQ��O�������$�~^,?�DPPm�YO<(��lJ�������A{t��; 'w����_]���;���;�ϔ'�����@ǻ|��/��ڔ����Β���kX��@����LƟ X���vCU`�7f6tE��e�~壖ղ0dr�8L���4�UR�����(3�Y�U7��
x���O�O�%q�;Tá���GvWOwH�j�N�X@�>��z��Ӄ���7ц���1eLڦ�3Bp!ȁ���'�.�A��?r��Oi���pI��BU˵���{<��FaCn�['3`vJj�(��-��������p���jX�gu���!N��)��/LI�t���|�j&��N�s��Z%B�t{n:���.ϴ�X7�U �0�,���,It�V�>pt��m��������ȵ�ml�]�)�6n���{{��@�A��r�i_���.P��f_����*ׅw+�5~3(5Fg�9���gh55���P1@#�`ɲ���aG!� ��PwD���MoC/+�Q^��n��hҎ���P�������aXb�?���R��"����A���,��ϳ+�6�����ȍX�SL]���r�!�O��?>�(ᄦ��L�E���`}���B��$"_�6�/�<�$�y� MQWS���8���9���7pi	����
MvZA��u���E�D���R�.�-�V�w�^��z�1n��C��B�AeJ�T<)S+sط6�1?�͍D�7�g�mgW��/���"!�����Т/�Z1��!���o[iI( iٴ��闐�E�&�j��^'ԼQ����b��� d��7fU(MA�u"m��b����K�G\B5��w�'�0[���cx?bW;&%���iwpWejC�]
B��\Y��$�6�4fT	�?@�	>`0ʶ�B����J<�;�����`1�${��X�T�D.4I��~͟eF���3��#|�hO���>��pq���wW�(���{������&��x/�	���#,������#v��Գ/DHJ�e|M8^����{��7�k^~D��bk_��.���O�5�  uQ�̛�P�D�H�@�V^V�x�&��F.��Ya�B���p����/��H:�򲿴���d���26��B"�?}u����kX���Ou�Hb�?K��;��A
`D���<6��z�I�"��H��UZ�y���M?K�L#ʖ����S��W��y��L	�ɕ�b�v�ye�ĕ�ǹOļv9��w3��"�MPny0ע������]�=��RE�ɼ����ys e�cF�Đ8�ط�:?��'���a�a��l���]�
a�1�g�4_�S��=�x3��b�QL�����ȁ����W���pId�C:GU[�Ѱ'� /{ѐ	��0����W	-5��3f(: �ͷ�0��=�<�-������K*3a��b��R�P�>�c�r}i�#�Q�4au�y�v�b�wS+��Bu+�Cj�3��]׌zR���5:����� $��$�8���+=�\�n��ȹ��/�@O"]b�ۻ`z�V[U@� ˊ���������	��s�+|��CH�xB��v)����YS@�,����9�?y�v����O��O�������X���:g�B����Q�~��j�8����kz�O�U�!p�Oo�H��ϏΩ��Ш�p]�r4��n�Q�qG��Z��M�s�(�_���4�b]�zt��H 
٭ő"X�XF����D�P�`��c����E��	c�z�dԠ�T}h��^��^V< Z�K������-����,����D���GZ���U�E����֣����F�<�����G���g����Y��7��h������Va��3��D���9���ۛ� Lm��'���Е�<��7׌��I�"�?�%�n]ˎ#;��m��FgL/��C�	�7.�֗�[kC����%�Rj�[t�M�k�������68.��%44��0��{ /�ZD��⾛2**�����e;~0/[QdC�oI#8/d�M��*��ز+��,�qt�Pڔ�� ��UYV���.�aK#ű��9J~s�0����;��»�	���T���fvl|Y�H�~���P�5]�����{l��K�r\��F�? �W���C=;&b��!H�Qf} �Ik#�PB��H�B���f/2��v�'t>1�No&�S9�s�PK7ӊ�	�O�DmO��l���<�+�O��@��>���P,ٖ����F���w���]���)e"O��\�3��x��iQ�����녻���\���x�|��ZHـ�y����Î�~��Y�}���������lLNV�,rY���}h��I�ۧ�W��j����D���?3aF5 Q�͈ �Q�la9�OӅ���Eۓ� Ƒ����y�Ot\]�6V�7�ԫ�G�oK�s7f�jl��ȜU���B�@��I�Rݿm��J��x�64Z���n<�I,�ay~�3 ��tmmy�*��:-��!�܏��x��0������Q�ѹ7��8�آi]�;}z(��x'ź�H�������/���^mT%��֖N����<̖ �6r�zYע�E���(��yR�h�?�bN��
~p:#ƳtU��ʃ$3���I��Z�Y�m�~�{��	����Z�8O���˭�+�m�Q���n��a�E�CWi�G�W��9�'���jb��T �1����V'�}L�}Pm�J*��,Bz.\-��EB4/���v����z0���`�*]�>���hG@UpEJ����s�1h�Fg��ɻBdS�:���+Ԯ���U�2�̕d[���ܱG�o���u��"�����ʢ�jߓOK�ݯ䙺�sG��T6~�n���tE[�l,�խ��$7�k1�g��Y�	0����'�I;�{�Vb�-�S~�aP�&��'��oЁq���<���@���4X�E@ ��-d`�\��R��w��������S�T4��v�����,Pa�d�*FV���4�����4hY��ǣ]�<��IA $�.��P+�"���i���r�Is"���@�%��To-G3q�����:�<����B�)�`�5�����#)�04�9T4��6�Fn+W%A�B^Z��W닚m;�K@�2�1�St������PZs�B�����_���A�K@�ȉϳ"���Y@��-ɦ��%[�`[���Z��B�k��bsg�����E��DR6.%:0!��2�<'�9)Y!�L؝�V5�Ǟ�!�����^\4�!�X��(�����nAP���E2�y}��O�dS5��eNŃ������)�&Nm[��s���e�P���n�-���u��A! �]����/8Q���/jEГ���EC?�_H*���0��·����K�<-I&Ɲ��ٞ�m�4�Lɐ���a`4/�2����2vF�^��fĄ��m�4E�?("����h���5� ]�7������>�NG%[�Gf�~�Mj�νI�;7�l�s��K��q�zt�;�uS��u�ji��H���b�H�����qC~���(N2�@��l/} =ET^G��U����<����
o��T�6H��<�!�y���LS��C$���e���҈i�D�$��~x�ՖiG�@9^k��p$#�X� �+�%�y�^e��0ڨ�>�b�ב�{DS���t��U�|]V��*���lG�<�'�Lb��A�e(��,�w�:�E(cX
�>,e�d�<�.r�����u۞�y�&�(CBr��{�FaT�]@��%�2Vv30��u����{��i�͘���G���^�wxr6y�k�+?�����u�֝
@ﺓ��C�|IQ��{�@��H���dÛ��b��Q#7�u0
�R�g�:���|��G��U�/6�g]�)�����xM�1�~f���ID��CNrc+�8z�ݖ���gY]�N)���''P�;�빮��Ul�c$ �޿������kpz4������8��I���/����l}��v���G.Ͷ���&c>��z���5��fs}R\j�x���O>�>���n��E8	�Ժ����n=թ�������*�ꑀB����_����,�"�+0�D�$�M�-bqa��)��?v�9��S|Q�aF����� ��j�\��=}��V��7|
�g��t�n��'$}���p���[V���Y`�2cD���e�9�2�� ș���D]�j�rO�g~�%)D��H[��R��Be�;-$h��K�
�J�����5���Y�)<�r�O�(��_�.J�K�󱚝�.��X̶ʤ���lǡ����T�}�5��،��	����rc��"6�{�$m͖��Po�\Rk��;˞�ƈBޕ*�RQ$���+�!��Z͚����s�m�LR@�T<a\��)�x����gG�8��z"�4m�Ǩu9�lK�܃�ł�
$��W�8�q�D�X�sX�0����I�.�ˈ9�����i�������a��i[	KW�5��Rj�,G9��@�E_��(}q$��
o I5\�ː9��)~��
��n�Zz'��V��,�Sh׸?�}�����Ӣ-|�e��L�k)���*��٧�[�L�3.�Q���N�.��&����ָ�=)q��E��F�#��^�?=�8�f�O��]��ob:܁���4�%�3���GA��&љ�ؾ��[y�h�� �������_��֮O�H������p��X�y��S6>Ai*��eJkX�ȈW��4�1u岮hķ�&�m�zDY�j�	
�O=(	!r<��e�����e���ԌA)��/!H9����C��J�|�A����l�7�b���'���#RgA ���~�d��	E0�&��*�"	/�u��]!,�w�v$��7���Z۶�dDӤ=��*1K���n����v)1�~�EV����;U�n(O���0�d����=G�8ec3{0q�����p0�C�]��D5�̔F��Ρ�Jc"y!.{MZ���{Dh�qZռ2�^_3��F$3�N�bi�V�.5��W*�N/~>m����wL�?�
��V�V~{����* YL�C��^�6}�H��)�T�X��B�Z�y����n�;��\��$�����ާc=ZT9��w�2C+j�A��xn�����HbйM~�|�/�,�5�-dG8dK���
;{�%��F��aw�rj�D�sIm���T�&#��}�*����m%��8m/q kwX�|&N��uW�����o�2�ϓ�ʃ�!hOͰ�0��"�4/qMǶjb��g�ʠ.�,N?K^�9�~"�	�(�rE&�"���d��ȳgd.�Cot��ȉ�O�9��H�5�J^L*a��V�+%���/_LEDXI���Q��5�M�tħ���� O��w)(�d,I����}Tۢ�$��I��$#OJ&_Waך�|O��t�����[�Z�(��T|�ϋ#vs���s<Ƿ�!�v����G����Q�N�I��,a���l�m��7����7��2n�m$X��M��gr���44�v->1�k���kJ��G��C��p{(ϖ>XPʻ��*ĕ.�[����Ԣ*�t�������;i5�/=���񒂅�E�RaN^�{O�y�
�����Pj����;X}�/F��B�T#� NA_�{�g��:�6Ф����v��q�υ�d������t"�5}l���h��/߿�i 髎�8��p:���o'�	�������ۺE�K�[j��5�N��|�;Q;��ʾ:�p��~ o4piUU��T|k+i�/\V�w�X�U���_�h\�=���J
�Rrut�0����'�苝T�.�TΤ06"���qr䖓�CAG�$9��(>A<�+a���!
�J'�~��8���[�U�7�Q�rC��]�J�r�+ǹ��s[�n���"oa�^e�B�`���b��Z���f#�z�˴i~nA�j�#�� �B�u�ݗ�P����[D�a��].�W+�b�o�z�UAz�N�(��Ն�b�O*��(��|�`���N�.�s������{�����*������o�w��_#kҚYt�ȑR9��[��K��{���8zd�%3��5�4��(u�>�$y�(+�7t� ln�X�~*��z;:��ͮq�C��H
�-DK;tU�'r��[��ݢN;jE�n/��:�V��W �]�̓�	}�`̔�<L���X�vs䙩!ѐ�-=+��j�o-�Pv�F���0�# \��<���I�}8޹Jx���7a�� ���i$G���ͅ
�G��i/)��s�:����Z��\n�3`v�b,�SE=.u	L8��S8���W��zs�j�}������(������@�%����ͯ_@�W��.�njr9z�wtպ�h%���v���ב�=��#ݶ�$k��g��$���y��ɶx�`�s�S6l��\����aAqW��z=�:J����Ow2	((}�)!;ʳ5�>ۛ."�5��?Hi�܆�g�����B�rש78��S�)?�a����=�>�7+�0X�;���Ɉف �Dk.Y,��񠄻@��:���~�.(�U:�P�4�Ӑړ���?z� ���"�r��9���l���j�әR����l�b��y���V~	ɦP�>���
3���\��
s�0�(�����4�n���5ߛ�1?�	�ֈEF'��V3���=`�4��ǫ7��]�E�4p'��gت7rP�!��H�F$�����@�]8L_����;�X�*X��URa5IZ�{�	q���?�;���q�:s��;!����,s��ۇ�3J}*�b��,��0x���c����=�*����?JSR��f͒+G�G�C��о�+T�`Y�#p,82L^�v�]v�YX^J`�x��% ��+$Cm"L��P��]e@&���-.-�SL����<F,��N�F �g������c�w��-.�Ӊ�>u<�8��G��.���#a�X���� *�B�����G��T����؉�Y>vNe�N�"�8A7*D$��#�ю�~&��{��4n-?[m�*<�5�hC�ѷ��4 �����t|�>��E�7��Yϐ��Tw���CN���)"k�O��7?�p���*�~W�ǩAE���3��庛�#[	�<��؛&�y���l\�%&�?rJխ@���۟tL�O��k7���O�,���N�z`[8����
�?��!��X �:s/FHϰ�������FE��{7�m�a�1wg�1�GQ�,:Wx�9���8}ב�=�W�u����_��^�^��Ț&�z�QY��ƌN��JU�LN��hH��=[�!�4���:L̺ �o	�.�9�;v?�����0^�~%��K�(�P*�ٯ !�t�V��KV�����+�uf�����gU��?CZ�a�F�=��H���4n�M�O���̩��i}��=�!U"�er+��i_���{oeQ|����8>s�Y=19d]����'ƬìJ�!� ��N��y�}RȡV��{x����� 3����^�����F]9
�1Z>0y'�7�`*h�j5���9�*��ܤno�Hk2�D0
~�xI��㹗fG��KK�]$*r���c�yW��݈"6��g+{������{ݍ)����es��۳�|�d M�-6��. uMl5!�э����g�t(��Z����doH7��LC`G5v_�3�v8���wDN�����������9x��ae�х)nW;�Ѷ,1�YH�v �,Xk���|�;�-)�r�(8qi]���� M���=��`Ȉ��(h@�6�iߑ1�
7v_s�	��b/�]	��'�h�o�Xi���w��t͕�`�q��wc��w�q�1j/�N@՗Cy:��eR���!����"qv�Y7NM�xMgI��(5���^V�Ӎ&.��؇sq��W�Ab�E�5,����Ϩ=���8W��P���w��x�3�"�T!�$!��h!:�gY'
�j����������q\2��/���.5�6K�C��[p;������ �M�s(t�Uc�����:\9�s��,�X/�J�e=�+SHnv`�T	��ki?�81<�2hFʣ�V�z���p��^g��G�5��D�{H�!H��m���r}p-�[xv�"����к�-���y�XuM�� ϔ�3(r��A�ǅ��8Xr�?}?:�Ͳ�Ɗ�k��9PJES��Z��K��&X�8�'��5Mȅ�~F:�&|����ү���s�H��
/��H�89����0$׀�`�`�XGk��T��g
x��#O�Fk�6����#jB̭wB�j0O �Ɖ%�^����8�i,cѤ����:Vu�q˺F�#��2���t�� tۦ)�q�N�,�MK����k(-�k�皞y.O^�
,;%iˡ�CK��i���Q��/�&����{W|�{��h���f���ؿ0�D�)	�6��6��3�đ�+��^�$3���$��oa�(c
��_n�r5쌝qIT�ӲZ�3���&�e��	&K�D��8&|G�=$��HAi?�a}f|umr]���Pnh?�M�&����yfo�Vg�.��J��2���O���o��*���c�}��NAo#���B�\E����}葝��MU��δ����R�el�A��uEP����>[
=��2������?�S8�E㋨�"�G���}��J���k�(��;�`>��IUن�%�ؤ�gZ��M��{��MK헿U^I�4�夥��M���Vl^���U��綊-ʑi�1�T�ї	��F���2�Z�z�}Z8a0p0�Έ
a�7�{t�Υ�/��n�,W~��ǌ@~�h�MѣA���<������ܟj��y�6/�B��c��o|#KTy	���µY�G��O� �7o�g��@�ĭ�o�6��GP"u�9(�+��#Z�*���Z��Y�ܝr�b�Q�w/ےNPÕ�l1�qLUM8 }��)����dsL�/��8w�R?Z���_\l��3���[��>�I�Gc�r=RE�E�ӷ/�@#:��'�\�^|A�	v�`�L��3w�YE �@�uThK:�)���=k��y_���*������:p����������о��6�\�5>H��~�d���~�B���UNznw����jb��V>\
{�T���Z�}�x���4@�;��eE�w"1�I���l�.S��J`���x��_GF�n�v*��Y��UĠ��2�K3�
w��]"���3�i�^���a��V,;�N���4��"��}DUGd����}/���ֈ�����45p��G���uÔv�o61�U�����  �:a���4��q��>VQ����S�ͪ�|Ќ5LuV����_\�6���>xU¨Oj3�Q�5�.i���u籢<NT:˯]�`
�+3�$|���p�>�U �u�Jȋ��7�����'<(�V�L��!�]�]nn�����Cs����){�B���	Ȏ�|aJ��j^2]�_��xxT�����.��z��p��Pt�Ҳ�.�z\�u#��ꀝ�<����G�1�-;��e�s��"�UBe���u�Y����{�<?�1�:3�\��%�1XԠj��+&��!��������Ʃ�E,���U����.��┼_p�AXerdY����M ?u�j��0�Mv]ZuAT�qރ�h�H1�܉�}Cb5�0R��Yv��H�� ���4��gb��A�������ڶiz�5#8������X����p�e�M�,[�:�Ƙ��Db�����j$��y�	aR�VC$�q��Y��sװ�耣Qn_C�P�(~6xQ��yR��=�-�q�U`����S�$�Ӣ�:��GHx =��ɂ²G�q����%	6���跬��o{��C���G�n��z���'e ��1g����ǧ�֫ڣͰ�v��BU���"
�����h8�#�J�p`jk#����%JPϗN�������#.��0��H]/���8b)Т�osx�S����7"R�����޵5�#Vw��1�}x59Z0J�e��o^�>p���Qi�k�A�����vIbhf�;q�����T�t�暁*������,��lhL��6r��7�p�ӄ^*��ձ��[4��i1��`�sJ>�)Vc�ʺ�?A����)�Aէ��)X�=<�_�w��SP1B�[LP$�iv�A�-W2X�L7W�x_i�B�C�����q�7+�����a�^ã�q�7�%է���x�W������b�|J�5����?azeVE���q#���Ŗ�T'8�\�a{�}H@����G�)��C��)+��Z���j�c���4C�b��|D����η�-��7��f�Y���p����7,?vÈy�?�֝��'|p]��;�ck�����:#�'�o\�Ԓ��A���_̱��VϑLܶ��˅�{��R��~s������V�@LEN{N0���a)U#j���gr]G)jh������[8�<���A۪�N�q���ܲ��r��������/l��8����"7ο�r������#�&��x�ސ?�d��Cj����S�u�p����{W�q��{�� �!?؁���m����#K�8�����+�0?��m+]�f�����呕,��W�(��k�<�e�f���:�������iM��9�&����@0�6��C2����I�6]�ʵ�����ŸĂٺ/��9K�u:CjRy�f���F`
�L`�M�p�m��oi��eN����P2g�v��\p�'m�a�,���vi�o2��/]���_�(�\M2QT�k$�#���6�wg�g��F_��*lˡ_fX��͖���F�;D�`r��y��G���܇�ں�{���R�m4.�%�|N�?���F̥%(q	��>��M�.E%,~m̬�${��nPA�U�=�L d�VSXH$�_�~W7��Bj����VM���6_�껮� �i�	 C�r�&�d��F�G�����,=�w�E�+�p��>z0P.�GՇ&F���
HЍ� Q
�>b=��pkz4ftA�w0�����{(O'k+�A_�٬�����G�+�T�oQ�Įl�a��� ���\7�l�m.�1�7�/����7��W�'����[AV%�FB���	��|E��¶>7���Y���Ԇ���-+���]�d�*���d����X����w��Nzך��N6R�U̙�o�M쟆�g�,1����SRϰ�W��V����ri&4�9��b'>����U��vÒ���y���E��?8k���#d��M��3ح])�j�~)�?�+�k���/��E�X&���P�"��7�`��5�S�uu��k�M�u�~H�.��	B�s�B�����wu$�d`�F�n|/h�X���.�榶���˾���zP�I�iRnB�Gh�V�[i�� ] E�5}�$軛���xw�E_>�� ��p;�T�;y�a	,P:�I�נ�[ �qQ�c��nT%���#(���Vߡ�c�b�BA�#Q�n*�0Jp���ҽ�j,ks��za�����g��:�~8ASOM_FL�V�h�F rE��8��z-kgz�n� ��;(�G9ֵ�S_�|��ݦ���T�g������Z`1�gTYX�a�O_ᕵ���׸<�W4�Ϊy�V��M�aI��v�b�����V����?�����%�=I��ҭ�P�[���h
R@��ɒ�	N<��
1�bj�b�wR�-��U����	��[9�p:��=v&�ŦN`m��n�y�<ٟ?��%i�220����R[��-H��l�/I����_�}��w���#'��kǆ�U�P�Fc�����)���-x2#�%��R�y��c�&����'��In�!2?��Z�D���;I��%[4�j��c�C�o���x�e�]x�8Fv�PnM�Ԣ��EG�:�dx�@�Or7��q��^�|����9���1���2�Eg�3�;����O%��b�he l���4�+A^��iT����J�+@���	@��D�n0"��K��-�J���8��P�dİ`S/)��r���J�e���}��������\�t�i:��ݹ!�9��n�n�C�#�����f�}L�ɔ��g;꣭����:>�c̀�lՃ�<$硃�-2�F�n�Q`��r�o+��S���@K�.���&1�E�G��O�.�}���.<,:iow���RN^Z�2	��LSm�#V����~�TUQ��6 Xw{����|<��L
/�a��9hQN�]��9���v��,S��#��]�d�5'�0�O���� ���p�gaB2yh�+�'v�2j�ךPx7ą�F��Ni�$��۟�+�D�yw_�b���w��H`ŋ�9�6!yX�]�Ǧ��-��v�
��A������STx8>�Q��
�[�>��"�Mh#ԑ%�����ЁlB��.N�`����͝l*t�:]|��m���d��t6�jB��6�����DJ����3=O�����B-ȂՑ�]��PDP4�z��d������2U?�*�Ӆ��$�U�%��l.�-V�L�����(�Tk�ڛ�2k�-�eEXOZ�X�OI�,�q���~vj;��ѠP���vh��}���P�6�P�9�n�'�����d��<���9��,W�,��f7������@�85��ۧ�ېe�u	D��w$����m�"�h�pF���r^bv��1��1}�Ln+��eYU�j��n̂��2`p]����#�&m�T�9ά[\����z�r`��`�7�nLl��s����2MJ ���vb&�b!&�Q�%���`�mp��P�ԗX~���W�F��O�*�3<|��(ܒ��p�FZ/��g�3��3���	�^:r�����|sK�����b/��/a�H����d�nu7p�5�6��<��1��NW�.�j��Ŀ9�v��
xW�ݝљѝ���=l��_��K���23Y/$���w��Y}�-����lQq�p�%j��O+L2������ ����~x�_I�������#�J۫���q�"��۩jw2G{�R�� C��╎�T��,g�=O#-��0Ꙙ[����*�	ܧ�7��X}:d��i���U�a۪�88`�}������
_�h�b��K6#Ò3A��v��c�f޳��yS����>������6�b��0}����Ⴄ���@�U��	��E�t +��퉯Ɉ��ȟڄ�]��s5ս���T#�ݝ� ?����sf����N���1�|!]>L�Gjc\��F��n�e�m`|����r/M�@,����VA����eS�,��BJ[g�cj3]��k��g���bOA-�U�u���m�A���S_hxIL$�p
�X��ukOHe�:Q"�ب�a�w��%����A�7u�3|¢+��7Tzwp��p"��2�֙L6c*����j�\�+�6�z�oF� &�G����`�~+�t5�* c�P���W�T����W�̄+ʃ��)bGAc0y��;�ӓ�O��k�&Ʒ\0�@��F�+-�<��+j�t(� y9b��Pn��*���?EpŐ��i�u�7��F��g�*�Z��'������	[���Ȥ�VG�����A{��(!c�g����ߡ
��f�IlA|�z1��n���rV�Gfٚ,�( �u9:',�^����^�Q��菚���������㑤�G�9Ò�t�4\�+�1������*�6 ���Զ`��!��6� J��ƸB~)��`߮c9�q��]��G�_��'O�hK�i���LAG$�G����@�9����<G��5CeW�8��bUI��r(nY�-�"L��aY6��G!H&��/�&�ո�=k8���"4��ºœ�]�R���G����q}�y�6x,Ee[����7˵�Z��7�1�̠̭�"�	���SٴA��B����7��.-���U8�"~uӄ��s��?����"4WEjqa*8(�r����("5<}!(ӏǁ~1%�$�%���"+�0L���RǛ���г������U����f's�<��]�����a����)ʍ����ڀ��w��!^ ��	CS��GJП���Q�D�?���k͒����؎)�g��}޺�`� |5�e:<�c��09���^��;ZG�r�ŀ�j�Q������ �+{/t���O�IC�FVet%����ȌW�l�ܟ������wέ��	�z�.�7���(ReIu�mK��HY�J���oY � =A�7�)�������y���.J�szɾN��|o�ZW�x��l�&jt�Q�V�2�Z2>����Y�P@�K�i���WeQH�����``ʓ�D�rҠ���>oџ/��_E�=� U>Q�h&�s4��쮴�Cj�_us���Z����Ѡ���`v���� ��u��oa�ԩ�����
� ���_���_鏤�2�uֆ@� ��7��(*QQ�&����)Ya��.n�&`f��z]��O졣���a�%]A9g�W�қnب����)�r��(��2��8+M��IK�Ĝ?�B�֗-
��m��@ڬ��1�������7�)u�bbWU�F�$�W�K��s�p�?����eBK�F|Y��*��o,n�Ŗ
��x�0p#�/�H<,���=��be�qy^-ASVJ̌��9�u	u�z�������pm*k�WsVp����_H?�i��>�-�~�(�o��z�k	�i��5���TJ�ΣeS����Ƽakh���魯4=�/�>�l: �U���j)��`�	�p}�4��9Q�/�w\N�b>����������'�~�x��b�'����'�\!��Jm�6P;��%V�kS���4�[zؙZ��t���47��T
.��ņЎ�
fPu.5?,B��r_�_�:��]C*Ƙ��Q]�6���B���@#i�i�u���ukI戠1,(�m���ؑ�{�����O ��D_g����{�>�&/ڭ��txJ���A���;&��1���!]�KT�>(��{�M
�XJM%�4с�Rh��hV#F��v��^�Al�2mp��G@HE�H(�1����84���?BV]�LV�K7�4�8Q���˱�e"��?1��%n�ۿ�X@靀	E.��KE���tx�
-���>ֽP[�<N���gg��RJ�K]NZ^Geք��]��}�<>h|'�Stvd;�Ƣ��H�n�_gT
��*���`X��G���Wd`A�5��ڙ���BѦ�Z�O�x�XA�"�m����5��J�A��rL̪�����z˞�c���}$ˆyٰ�����:������fl�fu�|�H"�/d�[�N@!T�}�����]%(��髳�]�T�0q�R��A8`�-5�j7�5���DUiꕤ�C�sZ<j�/;J�#bW��;�U�����k����`ҲK�|x|�jl��|�X�_���_C�W��*�8�UX���m��A�|u.�n�\��Q��׏ggp!������e�}��ЋM��,�y�1Ld��4|\�4,�����#i��r�T��%6l ���ֽv���f���ܸ�CG=������h<����^����nguYN�D���w`^1�׹YMd�������ng�kS3�y?`���֝պ����p��;�Ҵ|��$Y�l��^$�G�4��9���'$j�>eU�7��'�*����1�����Vu!K��L�9�_3�-8�'��1�^�p`�ɛp��ʳ�d���AL�5�M�b��/!ą~Bx�!>	���-���w��7���͓�M=��Y�-䠛w�]�h���#�Ų"}�k=�=�����cA����Ӥ��S�!E�Y�ZҾ�x��ҧ-�t��@~b.�H�h���h�<h�X>��V�հ�Z�(�)kݚ&���?�N�SS���?e��+*}�MtQ2���TOELS ��k��_Um ���p?��|�K�8�&Y7h��,�V�FV$>-��J6�ԝ�cq�
�)0�PQ���Pm*�IG����� ���{:���MW�ei��(�s��L�N`OA�� vq8�[h�E*��#z�UNw���2RW;}[5��7+ۻ԰�4E9�.�Q�����E��%b�W�*�2��;:~��M�t��4A�F�sCp4��
�\I�
���C��M�
���\���N�G3��^'r�����:\~:d���;��1�Zt�N�5F���fI��
�}�a�c�^O�浨|Z�lM����6y��~�"v��bճ�'��K�p���0e�<�C¨��ȒQϊ'
a�%j���lUU�ሔ�'���@�?��ɾ \Q`����3&�yg�%9���ZuwCw۰S�kJ$�+����).�i�^�pa�c5.���࿏��n$�O{���_��͖�n�<���Wqq�r|iU y��b�>�A�djN8b0Z�("tY�<��
m��1��?H�����#�=������Lq�q�h�Y���?k�D&��8��T����?�
Pq����U�S����� ��r{�$�s�ֻ9�D>p��s�atK4UG�&)|T���o�I?rv�B��O��hߠ��,�ߤ*%w=m>F|��	[e�Smn.�>̏h���̀C��M��YO�هTt��q�U}��OS��}�	Y	i�ˣAc��cy1l� A7$C/��=
&��Q��8�v��P��i���o�T�<r�!o�,=l�c�e�us�7�ʖ���S��1��^Φ�����h,UjS��aW���*w��%R-0Qw���xi+������qM��O�v�1GZ�B�����ѭ�9�����2YMo��NI�����wi��&�2a'SU1m.!h���eFhRѪf5�,o�B	���W��;]�P��Z3����/O�r�!|���E#������p���k8{���`d�^�H ��p||��w)�9��gUމ��ˉn]O�p�w=ψ=�^�r�Jc��Η�+���T��ח�K�+� �@���|������_����ƨ��i���8֞0;n ��@��A@~A������;�'�>������h{|ޛL�ԉ�$�r�S��>=���
�n��1�[��-�$�i��Y|( ����=������Nj���YZ���SyM�'w`�|_U18��9�9b#^q����_\�]+�n�ᗫ_��sͺv�D����<�j����#)��W$�K��xBd�M-/	+�>0�݅�M�
"�<⯚LoJ�6-��� �q$���e��x���PɐN3����9	���*	�$���m0pQ���P�j��e?�����wFEC���}M(�]��Ӟ�5u9b>�l�̞��*L@S�06�n�Z��L�6�0�)��M �Ð�΀�1f�a1�}��SFT�bXA�ɷ�=.�'�I
>	�|V�P���W���jM�����sL�V3�mH��kS�	��b�⸹�SI��SB|*ՇC2)�@���\Bl�7C�u���#�	 qp)�<��fE �e����C� �΋Lf�?Xg��0�N���%�:w�s�R,*�_��P�����n���O�m�,s��W���{Rg�k2q���� Q\���T1��e�W�����y��8#�2�ry'R�����l�������=��E~<G�lCO����9�6v5Z:^s�(�i��O"d�ƅ����N��&O��.P��ơ�mV�.�H�n�Q�
�pm�w���lN:^�������f��g�:Q8��3���)\E���6�J�<�*���e�\-��#��:X-nV�oi��� M�v+�(i����R���2f���2x�Cg�}�ڧ�x�MGәӋ�ָ�%?A;�m3��S�(�v��e��c׸X(6�ǑPa>�M��t׵Y�Jht��:�b�qWA Q��],9X?Y��GYK��j�Lh�E(�tzO���4�!b�3�|^��=V��j��Q�[�A�_,�����_X�>�p�pQ�Q���t��m���";�n��ޜt.U�i�3t#�@����t7~7d�!*��r}��� ԏ�;n��A�FS2i-aW��t!B�c����"M����D׍T&���^����d��%?�͂+�#��?�(rp���9�,f���>Z�������l��9�����#��������q����&t�h�Aȣ.����kkt��}���.���#��!�eue�ٹoH����Kz�$p_�}��
���0\�^_���-��b:��Y%0;ξ���_�j�~z���P����f�J�ۍ�9/�8�f%���z�Re�YE��"�r�F����Cß���>�9����"}w�C��m�T���)x��mh�fuyo�	)a�c9Y��#N5&������׷�������τ��H�8��� ��&s;�{���L/�0�,���#������I�a|�w$?�Ն�bc�����	�u;w�U���i�#��/�:1y�f�zJ�r��	�ϼO��#��_�19.g�k!�z�2��#���s�xІ'����Ƞ�ʫ(���4
�,���nAd��o'y[uu���r��\�6�x���n4����5̚�4ep�����T�N�� ��6�֥��˲3e�i�Z���S�t�71l��`���Dmau.cP�Z�����?��D�y`�E�g�R�6}���c�Q�U�]NpP���[����u��5,;��!��z���j�/@�����y���T��*�2����̆lL���n��0c7���x*O�
feGU7�B�G^b���Rfv�Zt1@����H����q�HÁT����5s(Uw�/q:���v��E	�2�1w}ɍ� H�u�����HB�<_]0eec��29��;7`����ل�R�iV���m>E�+� (i����hM��cI�����1�8���Kf9��s��O�x��b��	����6����̓�-�71��H�_��q��I�#F-�C��]�r�b��a�(WZ���y%O�y��m)��9� ~4��«��S����+�������+���m���X4c����� PD{�Qc+�~��3K.Ǌ�d�A�����<���X>@!��O����U�Y�b��~��� �KGˆ�¡�$��h���C%7H��m��V���
TSh6�*o|�����&����%A�Z�j�p' �-W�H� s�̄1��c:Ҁ�"�
�Žm{3{�O�b{�l���v�ל�޿�,�`�MӎmX�� 5��4�u�
�W�4���@���22*�!���R�'5���`����w՚��/��S�:����{�����bHCݰ
;ǻ�C�����`-{����,(����[��N�	��{�W�R+�������8q�T����r�o&hG�}9��-�w�Hy�Zټ<�ّ��<����M�St��[F�0��\����Ԛ����(}xGy��<��7_�W���k�V��9��
�r�fV�ku�9�d1wC�V
�}���ғ�1`,,f��` ��%���g(�^=��<�
J�}D����߁#I��W_'J��ȎӺ!�-�Qeo`A��6n}�1���G�������g$��L��n�X��=�h�^�tgӲ{]��@�ԏPb��m�X��H��s�HurR>Y��a���oɥ���3bW�0��Q`�G�#�e��S�7#�/UbwFÀ`�m�ּ��sԳ�pN��
�?�QO[Kri9ko������$�&��y$��ݝ�e��꛽�qOȢw8�|�/�~'�Ȁe{.Ӱu�%�]ע���L�h>��c�l�6�����]u+��4/ȝq��v��YJ���\ �� �1�9��b���v�2�ed�h3�=J�[ͲR�%�h#�|&��������{�:7I����b���&��s1��ل�i�#��	�.��6��Q
Zy�v]gL�/��Q���#�M���QƄ�T��T�IP1U	�E<5��"����a�(U
<f�����f�By��Y'�l�8kn����.ÓW���8��7*�aj�&oa%{s���W͎j-K�F�[�LV����+ l�X�4#�j^���չ��z�r�e�����&<Rm�%������,�G��C���X��qo0�~2g�5:?(�E�<�i�ݰ�Cm���ٍ��6 ���ސ[��L�{E*���#�v=_�@�$�b%����b�;��%�:���U���(�AN`/�"i ���mxs	ٝg��9{K-���Q�<��W�S��7�a�_&��=ws[�S
���a^��Нr�����=���C���J�t����S����ב-H�mFkv?_��iѡ"K �Z]�
���ɜo,c�-�Z	��
�Ԭ�A��&!�A��X*.C��j�zJ�����~$"�����������"S�^ڕ-�5�/PK��%���n�w�j�3�<H-�2���kw�r�:ƚ���`>�P>�E���j5`1 Q
��3�`���o���C�LQE�� ����s�BO��aΛ_�X���S�Fs0^�vT�� �|��}�ʙFJ6��=��O����1����,H�e��u�Rt��k(%���p�)#�pTl���m�L�̣$�Υ��t�h���>�s���A�#���<�Zq��Y39�����23�OW���!�I�L(��-T��
S0}�2�g�}����6��C0K�seO��L��P�r��T����EBgG(�8���k�m��7�C��6*q��b�C�Qp`�QB�>?\�R�ᕖy�����ϝ|��3讛L�Q�������=�o�4�$�����!�<������e�8�+0�3}������������G��L�<l�͡��/�ъb�Y&Ne���l���L:!7ߤ�.��/p��I��Jx�FMR����6�k����zQ�f�(s�T N�y%�9$��]�=�%��?m�� (��@p?�zg�x2�	�8ڵ���#����r��.��^��q1D��	�*��,�Xt���Zk��!)��Ӧ�}�99�eop�����,2h�z�gϹ������D=��1�����$Wl?�]F;��Ҥ��~�1�<d�Ӣ|Vc�ڷ�y�8�q�0�Θ�)�47�aCf�@CC��B�F�0�^󺂾/��-TM�~�%O�:��]�h����jt�(}�q>f��wY����G3��]pI�,O&��2������:J��
����g���tYW,ߪ2���|w|�2y��t����ʏI�i:W�'K���v���y�0�{M�J.s/$Ĕ���� �I��s
�[�`Q�y�f��ʄ~�y�s��}��!w��v�(����S�T3 nHJ��W��o���Y%�U��J��l��ƻ��s�I�񛴧��O<q?����/-�@�d!����2�0���|n��~���k`ԗ��y�O��n�&�J�v���K�
K��80q:���F���`���_����:ثч�y�}���m�#´�|�������!��O/g�rj�H�,�z6�Κp�����NɌ�ڬ�<8t���I���;�.�j�r����*�"�A�%�܉���ӬIT՟���ї� ���h9k@����%j
�Xb�0�,X��L�����b�n׈�2��Y�	f�r-�l��՘�ە��0�Jy��0���3�p�'��_�1�X�G���T��4
we?L�	��r��|����Ӝ��U����Ĳ1��Nf�ƍX���Z���y�y�7\�o��-�k �o��
��P\��o_�����9#5�|�T�_gS�8������a�k|� H$'YV�tj�_���Ti$q�^3N�������#p �����Q�d�)�;O�1�R�t�M��bKԱb<8m��}/�[� �/�0������F�����5=<�or7���;�^���a�+켁���r�(��L�)��m�q�b{����{�`��]OM��##�VA+$�V�u.�Q������I�tn��O�Ew��Jd�0|
۫�~c��u���3�_�C�"T<�WO�H����?BB��Hd���E+,�<�f$�J	���ȕ��t������s�(?��^Px2j�SD�Կ��4tg��jl�C���T��v.�MfH���@r7T�� ����9��$�D�'1J�������;ĬK&/ơ���| _�];{�͟U���c��{�j�矰�)v.̢!�<j�pX� ջD�ؿ:����YV�´��E_gܜ���4�u��nZg����+(p�iD�a��b"�xYR���$@�������cs���cd���ȑ�;� P����&�-��,YhB�Z�gBx3�K�e�Wg����`����[�$'{���V�x:����[=���N�j�u�
���ट�$}�,���]KL��O�jI��wf9�H���*a���Ȑ��d%��B��.@�$�2I<ܺ�y<�x�O��q��4|W.JFq��o6/�,�YX��p�@��k*�'�8)�;5���ҳζHk�G��qL{ ߅�Z��*?R&�+�ýr1	�.9�Z㳉xxe�:8j�����UDk]�ӕڻN��}�nWq�����ʾz��2y��y���stߡء��f�����6��]�`mZ��+��v�
N3W�;��!?*6���v�� ��nɝA�e��J�߁��b�(M�6��nY�SG61�r�.O{k����7>�O��J��d(%:�.Sc�͌�H�?MB]�)dQ�����\MF�b�;ϕ�^>�zz�?���SC�!3<�J&��_Կ�-LZua\r�媶D���2��Fh��$�X�~��r� |4�\�4��cH�?Z�q:��֒�!f�>�:���;ZzA��9�-\:&=���R[S�IxAx� �[��tq��L/s��Sx����)�Su/1��!���{�zL�v�y�X�mC�[�)��5px�Am��\�|�h=�[���t�;�m��<�ZA+Ƞ����B�Ɍ�%n���L�0�BŨ�����:���W8Ü�Т�ϱ����ʟ��t�S�!Д�|��-G5���!�L��:3,�T»��ǐ4����b��'={52���F�Ze���D�³o��8�{�a�%6t�.|p�wW]Gu�Y�J��������B�`i��CB��i��(�~�OA4���D�&5	.B�cR��g�Q�K���O�U^SYZ9�Qxh��OTw4f�ތ�h500�z��A���d�6�9�z*y��l=�˓M�}/�T�s%z9d_!`ƬFXZDޗ�Q]��[�t�D������nyn/jC�Ⱦ<2�={��ڀ�ʿ���R��4�sE���[X�g-
��O�ߤ�� _؛1X��t�p/�Z�\:R�o]�yA�z�Bm��
�*a�,P7X�Dh�ዶ��+4�W�=k���,����F�CI������!���Gy�Yb����Z|5�[�����ÈK�B(D9���.���@T��i�w����`��-Ƙp�&\�9I��X"�*�����A�ٴ6qlL�'��;����l�V�rεgnxm��=��ln�7��`�a��R~>e�RǠ�񶝘�#$e���L�
k�Y���p�#��|s�un�q���fHy%F.	ݬ��!��z����r�X�Kv��K{ֱȖZW���X�@}Ǒ�ӓ�|�u~ܑ�<�����5��N�|��6� _x���8�m 
����Ѡ!�5�4�$�#P��M��y���3��k�Ĥ��:lm�;K���-8��k�:߯�7��e81�f��k>�M�8dh���^��jW����u	�[q���e�;59)(o+[��O�H2W�l~P��:b:x�ӳS�\�C�/�$�rH-���&B�ޑ����vY���7'�PL��$��ڍ��4�孬�����n�e�1��~p�OEj�w?��	����6���[�-�����)�}�b��ę�sOl��~8����=��<�22����r�Qx��;{��v򌍲�bna� �
ۺ������ɸ
�����|�D�������7e�.	�� �5�����|t�.@>ef��J��Pg
L2nm������tQ���q.ȩ�@�W�)j\�K���vn�;=j��=�T=X��zN�-t��erE~ Mя�[�hf)%R78�-������^��U��������Ҋ12�8d7N*�V9��ܚk#�x�p�v���w#�y~,w-�������{�i�}�j���?�Rhq#��ĩ8���������sm{x�V�}8��B���s����x�q �~@�%j�D$�GƇU�cZ�fm[�2d�������J\���.V6P5�M�~!����5G#i�Q����,P5|᥯7�+P�7y�Y����q8��ݸ;�P�����=ʙ*��p�� �ܭ��~Tw��B�)�S�;j��YK�a�8�wgi��ZAE��;�M^�ԅp��
,U��M�Ֆ,�L���P����-ݗ�<&/�8ݕ���t�<��N쳬!�\�C�>2�q zmऱ
�h4��p��@/�1��2U�+DF҇�Sv���^����ːq$0'htn��0�5�M���̝.�,�P�8��N�c�1N%���������̺Ok��1��0C꿉5qs�(r�pF�(���U�˵�-a+c~ ��k�So�߸��?u���-e�&O���U�*����^��� �O,Y���(�Z�߈�^
�Z�����9�o���2�C�E�aP�n-��|��YR���m~�(x��+�UZf�׮byi'`�v�<�|�9�e^��D��9��+p���4k���s�9G#߭�P=�S���3⥰����طFMa ��V�V���q�Q�'pT���WH���L���`k�mh�����%u�}�5����)h��1Y�!z@����^0�c�tIa4���]ζ���89q�
���x+YXB�_)6��@bS��� e!,G��EVΎ��TDF��+.�;d���5��H}#w.`Uמڳ5��_^�^�܍ ?)�w�xXٖ0����Ϲ�ǮFQ�T�6<����%{��v���{?�݉��8}���|�,��N}mK|���ֶ?��W�R=�5}�J�jÿ/:��5�L��\Tn��+�z���06_�5���+�֭��V$��R�R�:��&$a������.�=��Ɣ�RT���l>G�ڒ���W'��w��%o��Ԃ�a�s4߿5���(LV�Dl�?����oeL�a+9�,����To�b��<5����m
2��K�u�23�����DL�����A,|�Y~*p�tT�(aɬ��Z�,7w�Zg�@���`���K�X�ݛ�R�D�קּ�r��k��I[�3�@�0�z�P_�U��@
l���8�E�5����}76O�Jc��$e�������b��M��s�MT�D�|G�ej�3dPG*^�c� k m��M_ŏv�hn�F/�m��(o�.<��oE<�0)�\λ���R�����w��O@%��6u�;g��r0�z�4�M��C��9��Ɣ�����ϩ����D��F�J��&	x�ui2�����O!c�SoFb�Z��'�����hs�`O� 3=��'�Y�a2D����SG m�)��~M%n"�l��{tۜ2�;��י��������Pޠn��D.Xi���܉�����e�ɳ��Cjs�	�˘v��W��)�x�9%要�#��AW�9�	v�Z������e�[�5/���+���?�����Hȩ�#`�:E���ƴ��!"�����#��S��X�I�,"�n�=wZ�r��^�)��%5��}�:��ʳ�ڐM��EW�z
�zÓ�E�O�!�����4(�Q��JUX��_\̸r_<@�G-4�|�<�6P��˧ҹ��G�glî�+�~�̷[m�[cg�R��6����0�߿�z$MX�ktҲn��@�G5g�V���7���*�)2�1	O��ҝ�a����}@]�����RW.IQ��	;�H���S��9��_�'��4�]�g'�y�Fh�������P��G/�"������p�M]c�ތG����L��P��st�,mr��� ��Qt]!�z�+ڗs8�x�������sR�Tt¯E?1�/o`�M������54_��ԯ�F1^U&k���K+A�x��^�q6�@��ǒ""|��l��2�Fi�<
*��b��I�1��7r�,�٨=c���g�w�{$�3ֹ�n��|)�0�s#�����%%-�yiP��o�U`d��4��d��5ؤ�h�a-u������
�F�����'��z�E k��膥�sjs���[�QZB�h�����n�7Ҭ�����Wn�31?>`>ͭ���9i`9[��Ა��u�3����fz�NA۽F,�CPDFhS�߷O�(-�b��mռ6����=�����mghܓc��>���	�������.F$���U/��F�j,	�%�Q����>�t'0���5\�_�oGr����?�}ia|�Ǌ;^���\�M��⿂����tR���CǦH�v���n[@� ���a����V��#�zʊz��r�̑<�K�4��\e�� )���U�e�)**���}���{�:���6�II1�Z�<��ȍ@�xK�0�)62�Lu�a��%~��T5a��5���`taj�����K������v�kv����W���D�/�?��LPS֚���C�`A��"I�r��6 %==B	R��Q]2u�}rR�4,fH'֘�a\ޏMNpuE���~��٩s����y��j6O��D�;R���X�� 0v�3���,Œ���z#��׷3#v@�dAs�c�*dI�o�u����	z/ �]�^�t	�::@����}��Q��Z^���z�)�EA4%�G����w�-=�G����*���L67�5|�iZw�<�Űh����5F9��f�k��@ƕ��p̚��܉�S�iD����"O]�������Ɉ�E����Na���OG\۬�wu/`�9��Cj�m�f�Ķ��hѻ؂��<��ڲD� 3&��;>�c�;�@�oV���0%y�/k�f
�Yh?���3�ZNW��ml6F�`B91.�f�+2���J&���z�(���P�%e�_ v�$��[��Gv���� g���J/��R�K4�i�j�Z�BJ�'Q��(u~��!)�߁�/�L���}��j����d}���C�z�����r���ZnnL����;��mώ�_�M������+��M��)����An@�<��\*�N����|�O�m �ޑ��hV"X;C��3]�H�	�\�3��g���*�5�	G���1̳f�ż�T���@v���=�7K>&ʅ�I^Y:P�ĕu��O�����
��5�X��,s��`;w�"�l6�Igrp�x�9봩-URAbv��b!�4-���_gTy؜Z��}=Pv�S;V�	 ?\"<�.�M?�vuXj9����b$��"*��ED�<RU���ģ9ytu��'4�`rv��
�sh�\�bg,a�w���8�m {��2
��'�H4b1����j��H0C�������j�1~�؊�;۳��#U��
c*8�-�/�L�N�ʋ��XQǨR�22�	�U8��?W������f�p��$44�wh|%��pֹ��8a�c/^���;T[�ޮ+0ۄ4�����!��/�Q:2��I=	�7C�~O��F9��O���.�t�Z����:�ĸ�χf"�AS�v�#o����Ŕ}�(�Z)!�lD;���F�Y� 8T�:��IQ].����*%�̃VA�F�Jk{�¿�CU��_�gx�������͊x�1o��1���V����	h1�э��߬�ql>��<�=���,&���O�Mg�o����H�j���J���3�M'�<�Yu��S<��F����Xn���#
��D��:�a��h��eeb�F�/�d������k����2� l1��:j0^ei@�cr����Ɠ-1������p���^�,�����5`o��d}�+��^�0o�3��;��Zq�)h�{y�d��ܢ�n"mH��`V�]0�-Y��㜞UA����5�ԑғ�n׳Z,z�L��ĳ?tx�8�q/�zQػT:å���c����|2�q����Yb�oO�SE} �j`�}�s��j��[z↰Mq�cxމ�r)�L���/�d�w�h��c����/�8��k:HڙQI�m��z��\ �~.`�J���@�+s����X=܂�[���l��lP���׵q�L,�J;����v��+�&�Z�[��i[d9�}?�_���M>�Dm4���ھZ��cBL ��Y�o?Q���Ĳǌd��ݫb�>w����h�-ۑ�a�|� /��&<���y�A&K/V�!��<�D�����e�p�L{�����3&4O�8�I�
��eyh\j�k���:%�n��a���G5��=ќ���������0�[-|q�U�����0UD3�Lm_�˔ڲbևC�y�)�oH�Z(=U�.�ya��_�{����*��8�m�=.�,�Hkط�Q��3�ο�q���MTD{\$ �!��8�d ��~Z�I��,�����8bq��U�����z�JN�Z��k�wO&�fq��*K����8�pEn�@dﴑr���ޘ�2I3d,E�����J>���=�&|�x�ě��:ܮ2!��z�{�1=G�k�^[����LP=�3�p˜�e�h��,�=�$�G�Y�n9�l�0�3wTk;y��B����zϧж��,���b���Y�A;���bF���N#E#ڒ9+2t��Q�`M  ��������2�w������;������+QV=+�G���9�+�50����ή�:�}��?ɮby߽£��$N�k�4(w5!l�����Fۊ���5����K��d̍�p�$_�����d���,?i|֤k�l�����1ɥ=�y?!�����I�	s�d�����s���+��[LkѢ������뜢�+�|���k�_E�"D��`U��b�5������C�՗я|"G|k����Y�FxhMr3v��:�a1�����C�~WS�&�&��)N��d�Eg9�X)�f�ZA��#w���,ѹ��W��s	Ծ����GH�o���f��I�@��3���'e���=m�k�9,Ϣ$��39d��R�X�Y�1�!F��8k�:�1���(���۪��lo��`�d��*!NPn�+�H�]va�� �V��u�U"VVz���CaIa)��|ҙ�Y-��� �teD_�Y=��YPK����3�	�%[1�oB���"��L,3����*�v�$�u��ֿV���W[0^�gP
�WضG�9ӿ`��=�I����kم�f���Zrvͩ�M�"J���
&H��]��f���)�F��L�P!C���h\D~U��:IVR�P&�=�M�y��$�GV���0T��1���罰�勸�a�m�c6~\&�¨N�/�.Nti�_�R�Ī��4�W)L9��3iE�ѓh���$���K�|�C�����..�rŝPg�z����K` �殝%�|bE�b��,�0>�����4�ѹ��7���r�%@��:�t��D�"[Y&�c�ZqȎ�9��"mZ�.�_J/$G��'_K	�9��i�㫹��L��3_�<��q$(BHa��[�泯��v��� ��Ȍ���Tۄe�%]ե��FhO��v`�/�⯾�T/)�5i
�AVx��谉�����[�nJaXi%;r��9a��]\�����.¡��87U�8���3�	\�E8I����>�n���RY�V�Yv�`��C��� �ge���+�Bq<�����w�G+)&@$?��[A�{�e\+��-Cd��iEUl�^B���o���|l�p��60d��=z}2>S���J��'n&c	�!���ܠ�9$I��2�9K���7������7R�L�*G���&I�V�
�|����A���9�����^k��|��N{ڬe������0��X�n�P1w�� $O��@�%J:S����<��qd{�D7Y��ΉuJ�?�N	7���:��,���S����� �^�������%el�ʹ�+�F�/r��q;ի���b]Ld��+N���#j�;�<��bC	�{�6\*}�W�����������9bmX�BV�����QU-��:Bt�2q��fxi���[�Q����Q���JC<o��[f�<��lNOE��p�.������	�[F[�踧R��Q����	0r�#&��ƍ:O�#�Uw����1�؁;�PY7�LS����"N�O�ˇ3���
�Ȩ���:�<`V}א�_�����. T��0K������Iȑ�����{���P-�N�����Eds�ܷL�����!�UD}�
�2PwmC���h�@H��/�����%7�R˿"Ç�p�O��Q��g^d�M��ʥ���3D�Mh�<���p�ǴV"]j�_(��Y4��`x^�e<z��Z��cCN�X�!��L��1��Һ��9���I��~�g�>��k���E͊���I�V�9�P���隭�S���x&5�A��
q�����
7��a!w>4\9�Le���Ү�χ���eg'א(g�51�UQh���iQ(EG��&�%���)��[�k�@2��慥Ih<4�����Lj��C�*Z+ j�ܭ��9}Nްo�#$��d`D}+��n?M�I�wNR���@�o�K���m��r�I�C��h&ھ�_��e�	�d9�<�j	�����Y��{���Ē��ny�I�N��<;3�8wx_�����L׃��������$M�JY�<`]
��mɶ�4�T�e�LW�.��,�$�#��t~�	X�S(�L�u-p���2ivMCJ�8�0�ܒ�,����{�ZP�M���b���8?jP.�8�ISD�[�k�����v�ZA@��;L���6�t����|��=��E'K�"\ږʶA�����
a��-M z֞w���^_c
V�6+(q��[��k!��v�ZX��d�A<O�]�U o5mn����gN4S�	s��x���LA:+�.���c�g6� �T���Z� h#�Ξ'xO�ٖD�(�����¦m��� �؇=�3B��y�N�"Cς�'���u�N��N����[�Pl浓pu�(~���3�D�Y����&����~�xv���U�;���ȼ�	��+�T���*%O�;Խ�;�yeI��!�tC�[�O=J۲�0�*"�ؑKr�G����ϙ���a�vYd���m9�*���|`��gXl�k[^D_�3º��ݹ�P��
L۞�D!�?�m��u�Ҽ���#>C~	��ւ�E���є��^��Fڜ���e���,�!�
��4w��@y�kE�g�Y�Cˢ�R��N����ڙ'q�ٍ���7���%D��"�Q�b��O�7K��#���U�4幗�7�\*���&�q�ݼ�Z�������΄qi������{o�-ږ�}�εaC����a����:Rl�WܨT_z�����c�͹^ήؙ�� Ms��|�&[�UQn}�jg�ZC��Om� �DXڍ�����:DDB0�UZ,����<�������^�2"��;�����7����c@W:7����ꟀE�}t��I��	r\�����/���R)îހ3D�t5�B�V��bV$���쁯~��p!<@���1w� J0�T�呞]i��;��(z�-/,D9}D���WU3ӕ���"�0n��iG��WZ�IZ����zv>)H�?����\��u}Ɋ:fmF�]o�.r�Ԏ'��������`�7�a���{[�%��꼧R��/�c�7����(u&[2HE����ZY�*~��Xt��	�e'�]3�����=T%�?l�����8ׇ��m�9CF:�.��L�"��^[D(�&/9xY.����I�`�u1�y�/��bk��ʰ�x�Ol�l���h�:�������;h��-f,�Om���`{~�	ꘅU�#0}}�L�E-� pK����}��,~(�����E�x�k��U�N A��zABsŏAz����Y$˽���l��p�Z��~'��]z�U��К���*A	ZE���)���f�R��b��o�"$�֒.j�F$�c9���6�I6��ٳ�)@�fÂb���p�x��͉9��\t��0r�F���1��M��)��(����l��n�`�0��V��,�=��D���y�J��]�f�z��s���#sR 3N�� /y��
����{��� �������K���~��L֧��l퇌�	��i��?ˬ�r$L�'�N�Y�$�i��b��ԑ��N�5�/��k��a�Ѳ=�:����u�k�(j�j�-L��:]��8ʐ�Q�l��Lsn�Ã@<}�e;�3�D״��v��:�-�i�|P\X�������5M���q1������8�WmN�更27󛿅lЊn_�����r������>t������B�X��=���7V��R�$��m���n��v�}�����\a����2�ݫ�!2ql@��sBS˧�������"�1��X�1�#B�c�{l�O��+�Y*�L46Q�㮿�W-Efa�>6�I�(	��a�w.8�� ֨�-C̒���CH�ͳ�1e����1Gyo�BvQ�e<��b-]k��M��O3В�#$!)�a�Q��D����ꌸ=q�˲�1��e�3]J�������E��с6��J�+?-P��+�·����J�M���N��FA��I�һl�\\�\r�����@��(q�ar�i{��e�J�f6W.���C[Ё�ag3&eG�0p.0�x��9#�r�(%�$e%��gѿTlI�F�}KaB\��x�챶Q~�����£�����u���*���Y�w�v�=�%�+�!���<-���`�*�,��g�z��5)%}j�\v	��Q^Pq��7����)Y�&�0z+(D䯮����m�u��;��tI����~ ��0�uwB;=%Q1����2//�V#��2��3`�W���_�$�=����O�?�H`���H3�)�>`�6���b gT��_�X[L�~ƾ�[_�z�:��a9�O���Du�3ĳ�X#|��,,�Q�QC����l=TF��m)�1�6.��M�.CxC��X75���Kb��]����~�m�w0�?d2��:�Ќ� � �p�я@�O+_�.�����APD{r���A]��`hE&�d9��
.f��B(2r��[z	%����ܖmW��@��H��5����g;���Ɂ�����m��]���e���`�:���RgS^����&��Xk5��j?*�C��v��d
35jK0�j�+l�E�(�Kd��Vd�����R�n�����d"q~~���Q`$O'�)E���8{��������}�Oi��
;m>��c�����y5�1�y�{Qn:���YӐh� |d��^`���眼�kB����j|ھB	��ʹL0t8xvAM'H^0�9��94Q�*�)h�pgX�5�Q}!�]|"���u���C�H�\�@������sn�5vZVѷ"^����#MQ`�$� �Je����g����k`�ܕ�+�Y�@�'MX�X��)��$�Q�#��<�*��y�O�����,�M�����`/>�9�5C�"<�>aP4�A���dM22�9�3�j�/=�1�T"�+KE�7uy��#/T����-�Y��X=E�5Y�+ ��]�;����6Mz]m�H�e�܋,^JO�>�%������n.�� �oRm��n8th�22��X��W�q ��V����[�]�ou���3�������-4�Vy P2���
�Kjk�5ם~�J����*x�J��n�꽇�)�UבX^l���?h�5�G�Ӂb��� ����C�/DP�f8��"d%�����G�P��P��`*�ȷ�8yw!���ҍ�'o����,{(!$��ƊW�`�b�~ᨺߠ"���_���%W�DI��=�����i˞"��=&������#^���zf٨f@?I������Q��7�G~����2GC�r�7A�Ra))�s�`��ـ�F]"�y����{RFT^E۶���#��ʭ�L����wb��9�b��|8��9����I���u.�A�>��K��`�6k-��r�qR��k�Ak�l����&y�l_�KI`b����{_���ؙ�/�U.N�9�D|a9��X�p�4������BΣ[�'i:�8�5nl㹎/y��s �|ȣ:Lf&n�ۑ�Ԣ5����$�D��<+�[9[�+���h���:��N$/F�5��FA$��H��U;yn�������/}a�o3s���Ms���rb�dQ}GΧmM����p�e�Z��>�O��ve�>|�e�5��L�ǏǹΤJ�ѹ7�Q�8��R�g!]��B�=�U�����FPuk��#._2״��U2�)&9��"j������|n
����*c���S��>�pMn?	���)eu#�L�.�+]��ɻ=��� N�*o�����Հ� �3-G��-�{EP���Ԍ�$�� 3W�}�ݷ�U|P!lL	6m�s�!��N�����b�!1ǣa��؏u�P�u�R���1E��/�S���,��d|�S�5<�dDN�L�W�%�2%�R�V�L��I��fg.Z��ݭc�B?�
�U��e�*�=07��!LV>��\H�I��	ş ��n��ȩzq�چ����\)�w��4�e!$?�2G�5e;&M���Bw
�K	�w�`aH��©���5|�����anlAtv)Q
/$m�ɯ�h��ޱ�h�X;��R!��r	���2(���\P��s4���<(�x)	����9ˏ�,GRX�hf��M�K�Z��
�����8�|]�X����xF����?~���P����i} A���ŶW+�d�'�8ս�Z��������=y���K+�v�(5�OYt7�H�b����
T7�{øZ� l)F��ʪ�X����b�K&�!4{�HNx�t 
P��KGu�����o���4E%�4R�g��>[�suq��mֹ�`�VgO,���G?|y�/\㳝����d��cm�y�<�,mJJ s��`�B����0FEV��?Ҭ�M�v:�1���H��hx�ʂ��H�����V2~���F�H�|�;*�T�ڛӒ��,���
��7'cgk6|DOB�f�2�5s��ְ<��bHP���P�Zύ3��e	o� �	���K�y��uu�}��'|���!������	SK�9/ �ٮt 93�������©X����nҗ,u'����d�N����ȟ��u��~�5�䵥�ZRm�i��y�x'���2,�L����5��r)[0M�+L�m�Cf��<(S�]�ᖥ&�z��L��\4��?������!\��U��fW��v��2�Z�)txE"�sM?�r��?����G+N��]��B�'_���ep��(�")��}hE��Ք�m�����$\p{x���|^��`��նCo���+E?��b���J�W����Og�5&q��G�#��Fȸ?J��g��ժ́��֍��{�R/h|7�/1R�tQ�P�	��)`�Dܷ1H5�@;Ϗ0��zdd�	a�y4�_����t;C$�$R�L@�����1��L���i��i��(F���Vf�Rly`������?�VY��ͧ��ۯ���6[fӴ�!Nģ�	.l��x�wq9�CqMj@�-�}M'�9M,��������^�x�~�&K�l��
lmWF���8�����T��EFw����]���H��m��eA�l9S���Z|m�d�`?�e1�vB�K�c��1����߼2���ߗ�S���0�b��	�G�yURp��o@��O�[|WI�E �V~(��[%$*�f�l\�n�<��Qr�$j���%R1n-5�`�'< )5��B�=�wd�Y�6�����&n���(�p�FMo����f1JJ�F�S�W1�Ԛw4���04|�e�]ը���A6��])����H(� ��� �D��7[���^�(�R��qK�pØ��T�l%���C�].�J��l����a-��M�ջ�����ji� ��$��>hB'
��V%��A���ɯ][��6�@��r�G����l�!��C�q�fb�]�M_��mIM.��<^���(�s�����V�vO#"U3��������W��Ai�M�0t_����<e"��^,�'�R��w�ӧ^˘��!��3T�z_�x�qJ4�����6X���h��3u��ѩ%�	����j�s��T|�+%�����cnA:o��8j_�>Z����J�E��X��_�n�0 �m�$��Y��ߌ�c*eoW�����1��}���Q�Mi�B���z4��LJ����H�E5���+����?�a&���o��|�Y,����{�w��h-W��}d:~Y�(�6��"}A���$�D�D����w9!ݠ�(h�﬙�����>\�a�ROv���fj2/,}����,>g7��y3d�N�%�:!��>-���Z8�E�R��h'�1��	b��t�M��8��F$���n�H�{�$��mvV�/�>50dzD�"�*���~�(6+Ǚ=� #�̕k��r������sVj�)�[��\i��o2ҕ(����lۅz���� (v�B�7}R2 vcV��ƚ���<o�}�j�p����K�o�8]�)����}�Q-��3�z����^��d3�ۄ����Y������4���DK���O�0�b�<��Ũ�~��&_��zap#�C+�y��&�kfc�b���h?��_�tNV��ܒ��������f�5w	�ԴsL$�s�.����WQ��E��A�68�EqO�p��.*���j��N�J3φ3A�W6�Z�d�
^����W�Ϥcp�03��Y6�x����`h�>t$'�Y�ЛH����KD?͖Yy\�2�N�r��U���K��f�V�}nD�TdI���1�D�I�7xZߨ⿟�\O��4?��9����}Dy��.~'4S,9�ϚzD�J��OW!�7�����|�4^:7V�������{���*�裈�%�{,������Wnl;��q�7�]��ݲ,㦊sсWJN�f&��Ɉ��:VȮ�+�S�i(%�}�w���HF?�e���N��i�V��F#T�z/]�"��o���y��i�ٴ�`Kb�^�1����ʪB+�<(oB3G2`
Z�r鷔����w�D�8[*���C���)�6����S��X�)�n�l�'H�Dq�q�Q�`'q+CP�����AU~��}�/e�k�}2�e^��?�x�y��1��g��D�Os�)N��ӻ�����'F4�.N�>�
?;�_na�nY�D�|�c��kǣ� u�KQp\칖����SV���� 0ׅ\����q��k���}����:����op�F,�{�4����P	s4����jw뚓�ykB�z(C>W8��=��jX���ɟ���5-����AB�)���R��u���̬��������P�� ���2L����
ߛ��o{z'�n������hi�����t^��T�H��UCa�P��u`	��-�c���)Ɩ��2�_oDQ.uD�?K%��2��ct9n�c��]Wrk����o*��a�Fu1�|��D��2-%�7�Q�Q #�V�-W0I�u؝�����Z(�ȗ�+�>_G��2��A�Q�sԗ��Ϟ�[r����f�/+C�l�˔��j���!'��u�Z.`���W���P��ȪV^L�}(�����m�Tvdmop�B��L�wm|��9�2�_�� %Ek�!��p�R�vJ���6��fg����.��IL�Wp
W��B�:��<Wr)#�ZJxX8b�L��+���aL?��� ��ü��`�c��RƤH��ڏNu�{�����,�U.L�jf�+pi�������� �p� �Y��R� AMuZ����p�l�ڢ�߮��=F׉|I�')�t<$^� Rr'h�M���}�R�9�������?Z��G,�r��������)�:�$���1�CC���x�b\� .�0�@�1�m���
���:e�����O��Ј��_�{O�璍�`k�}r��S�:�O����]|��J'zb�k
�$p��4L}��7���B�n,*����-k��X�"�rZ���\FYSp�K%Q}�����X�qЖ����� ���0��{��\�pjq���к]��$쒆��2�yFg�2;�96څ�(�=��//��~[��g��C�撱U �H;I*ai�_eP�~�ރlC�M9Z�s����$�J�Jҧg��%�S�����!DF�`<|/���,�{f8��p�C�"v;2��
q>�D����.<(�������Q��N�
3�3?�Pj	q�p���G�I�ܻ�h掀�T0�+� vH�#�t��7r�'�e!�R��j� A!�$�����rq�&�<��lu�y
�;�GV����,BJ�d3,j~����y�`��� *m~�+������:�H��MѷVz.�Q ���	��-��:��3��BiGi{��Kos�n�CD�]���akk�T���~�/;5G����w��g\��aa]L�s�ۄ\�ThV3u�b��楝�嶄��q�g`��B��c�"eS
Ыy�Js�ER��s0=��;�NH}��!�j�[�N���<=#,8�\1� ��ؿ�Ǳp��P���z��B㭿�a0r�*NW�h��a}+�����1�"��˳7F�O�!hR'�J�V�n�����!��R �2&34_�(�DQ��*��k|�5+;\�hMe8x��c>¾��o����Oh�ƾo��������\�7���l�m��#��px����q&>'�X)��S����,��>6	�1�$��l����y���V��	S٭����pn���=��Ҁ����3�!,����l�f0�ؗ	 ���)%к��[�� ���x�XH��ʎ2)\�"��m`���C�s��4���E�Zw���#A�sL�h�1��*W�[�J�&�SA1�S
�u�>�Z多c*�>�'�`�D|���`�h]�����o��셑���Ar�X��Wv��)�p�H��1��?��u0�� /�_�D�p��b�Nhu�G̬�Y���nQ*����A �\��*��v L�	��V.8�LU�ѡm�T���-j&����p_|���5\\�P�B�dB��&f����� [����2�S=R�8;�/�j���u�<�z�R�z��Xs��6�^-�"��ц
Ҙ�/;Uf�7|V����뗱��1�Zl
�o�o�6QU-09��T�jH�z��\|�A=t��.�c�JLV�.)�h���0~�5�0���%��z�:�@��.���, ��#}��^0#�"Eu��FȞI+bhV����cᵽ�A��;KT4��k?�o� �vEMj�pW�o��2Hr�FQ�JH_��X�S�M�$�l�$3e�/Qz��4K� ����yyu�sҁ]���zэJ�P)�5�� ���z� ��>?�ڸ �>bT���/ɋ�v��랢�/�z&��O4,��;RB�F:�]9�-��0�ӗ�z�91�e���@4AH�8�Uҭ*u_�!���dИ2���X��e9�k���D���f�s��ݶ�\�����J��#�P�N	�7dnW�㓘M(8�G�>1�S�M�A\���;4| ��dB(���������k��Y�ӿ��Q�q�E<�Kprq9.���:8�߆e��{L_ �$����E_���v���B՞R���(�z���=�Uh1?r��@y��Q��B�
��n�#��I�In*��n���������|����cǵְ݄��y{���}7m�W����i��ɿ�R����#�t�7Ɲq��
�xzIM%�PoZ}l����Y5�����>�]-�����o��bْ���WW\��d�ad!�%�Z�z��9#��2₍)z���>�V��)zBN<���F�ٿ1�p�:t�yo��o��>�,%���+p<�Z�c+���7?��1W����w�䩰l�`�Ay{H=���R��Ol$�X��x�[腋��NH�;щ��^͕\7Ld4eQ>��c�$=�����.�S��U���
lS��A�2A$��UO
�;P�g���r�U;�,g;�[d����@����|{��h|�Ɓ̂�c�^���GC����Ƿ�i�;C��x�9���^a�S����FN�W
c��*	&|�W?,W`s�,�J3s.
�+*�2��`���leceN�g.f�jʷO�4��a�y~͚�c�`�h�<�boW�\����k6��F��-�����������P�Q�WS��3�Ր�4��7��$�W��QQ| l-���%k��:�`��6��M�o�q�1���b_u�vM%���M�'��0]�?�T�30�3Č��n,)F{rs�n��'��NvZp���P{Y���݀8���r>��Y�����e�]����5��]i��d^e�g�t���L�����S�ؼe	Z�������7x�ˏ$������ԬK}U���Q����lF~QFV��hL�T6������-�&7��Ŵ��	1ԃ��0ӄd ��{���U]6l�B<�U��[x?�ڡ'�*-���N��+�����5�y�㓢���{�0W�*Hg&]d��e�� !G���2�@b>}i��|���K�,���o`�Kэ�m�����lP;��8W�4 泊�sz��k��i��Í\̮�h����n����\R.�qv�8�Qޘ��+dJ?`�S]K���ҰW(���l^�Y]�}-�N���O���L3s��9۴��2�����`��U� ��'���Yem ����6M����B�C��ZQZ��71�۱��׷�,'g�Pn�ǽ.�c$H�q��`�;o�0����o
�RW�.�©�o�m�5L�%�/v囋�3�$�!�I^������sbu`�U�|oǹ�	��I�W�����VʀZz$�����0�M�Z�'��>��sE�@��w�ƶߓ��2�Čle kĩD<��g���m�C�F�z���/A�T-M�ㄔB��d¸/�:"�xf���Hͻ+�G��9��?Ő�/��6j����2�ї\?^�7%�!A{w����(գO �R��E�����]�u��p�7`Ҳ&�O��9e��鈶R7{����s�7�W��;FL>���b9ل�T���m�z��x4�jV�"?�����ޣ�2�G}����m���D�D:t^YyQ1��?�����dx
����s�G��'�e2��������� !_����W`������:��V.�e�=���y���	銕Ow��1�WXjT��%�}o����$w��d��t	��]�ؑ ����$�jY�'F^Ʌ]�u�)��og�.9f��<�ʾ����d�x=��(J0u)�ǢS�̠�-��v���hs�ǆۼ�@-r�釺�3��������)��)Fh��6\�t|L����?D�o���U%Ϊ��x��G�Ͽ����O�������`�{j�lÆ��n[豝���dR2�}����0Ws�j�2��BH)�{�$ǘ�����v���T��atYp��v�S~^�2��[���t!�ȫ�U\R�?<>� ��=w�����`��
���z�j̀�G�9@��u2l�Ɇ`w%Uߣt�ߥY��7u��|��� �+\�}`���M���H6�>��hE_�q_�_1�5�)/�򈱤j���Q�>��u-���z���U6E;FjX[^
ү�T�*�j�����|��?i �J�:�5��!��K�8���ʺ���0_��LYӑ����iZ���ܴ,����T�t��]`�q�p0�-V ��}���X��q�JL�0�
��7/r6�rEO)5�(���ź�A�-$��XQ�o�������V�b��`���p��2�Ǻ0_9#Gn�g�E@���L��L�t211[���7r�)�LlQ`�]{�pg#��|�'A�3�<�?�I�I��m�M-(��}dDO��M���AGQ��RIv=I��ox��l��G��&������pԭ/ɕ�����%D�Lpav�ϥy����l�������5z�J{��(�;X� h8P��9���p2.�|�B�M�Xy&��g$J$�<>�]i��bS(H�/��9?8�%���L�O�^ۂub�v,�~q<��Y/��F眯%]��k%��O_�)�U�L��iS�B�:rK㲹��*ą6��T]�bH4��Ĩ�Q�u��I���a����eU:n����7X�W��$еޓ�4�����?�gJ���H��޶s�Jp�K�YBS�y��F����)Y���i�Y:'��f-^c����t+ /�5a�{��-�M��pWK�BSW�0��A~T]�dKz�c��a$Ȭ���T�a��9�EM�|gKA}�#�hq�-x�DZ��^�$@)m�>0%9s�w'�l����l	�X��9�U������6x���7§̍����t��p��yTpDi�#��+�]�Fbf?ƭVu���6�܇rQ:>RCٙu�n�7B_n$��ʣl�!Udq=�#�;!��q�&?S=aпw�\�k� x�@��'}{���=Cʨ9���.�6㐼���_�x֩�a���X�wn=����������XKΔ��V�?��C���eمCz��"S-G�o�YX�[��C*�5�#�rTZ���e���.�]a��	��*d�ʰ[�!(g�on���l3����Y����tm'�Lt� @U�ʴw��C#k�V�Q��n�8�8��ꨧ<��W9��J�w5
���@��+�#��5���}o{'���e�b���-�q2�#S�x�/z���x5r#:u0dO:�d_*o~\��O�E��,���	5Q�Rn�Vy��u˖tG�{"z���V��}CHj�J�<�_b�4\�@{��-N��)�z|��K���P���0�n�V�4'�m�\ �p3;a�/ʢ��~b�.����}���0�������|U	3sŗ��⪃R�[2��N.t��N",.�ne�%>�xN�i���uD��\7�0�Ǘ���S
� 5�/�����{��������U�����T�\^�h�y|`���J��m��Nr��ߊ��kc��W����h�`2�v'7+Q)��84]O1��/-|� 4��i���.�m�l��q^%�:���ԣ�6%>�Xؕ�3�;�<�!���ɳ��6HdM�ۑ� �/�*�zXKI�ъ7��G��u��Ҕ�g�!�����kU/���%�V��S���ײ�Us�����e������3�@:�N�O�j�!�g���7F�XS� F�Y�V7<��N%}@�WO」06�A�\X	Օ/-L~��1�۽~�u_WЙ��̘Jj�8l�A�#zʜmi�1j�@r"�<>��!~��@��`��0un�s����C�����eV]z�дk>jX�|!�؄2�{��$,�lbVKb�y�f_� �I(hh���P9\��c�1����
}�W~�\��nV�^gѱ�Pl Y\�pq�Wg�`�%l�`O5��=���,3�ŗӠW(G�����z��c�/Y���7�5�0N���s���<���mTx�1f��;x��G����9�����<ﴅ:(҇��fʣ�T�=^����{JiI���a����������ݽ������d%�³xl�6�����V ����^2?]F��E���P@1�Š��&$�C�	�)�,V�F]�}j;���k�URµ�!;�#w)����鉈�C�������/��w[Ԝ�D3q����\i�e>� [jsw��;)e:��u�a�b��YE8��9@�$�6�k��� �<��*.B;��̨���{�Ա��Q���!��Kja�l�/<��n#se��`�Ed��vqK�H�gSX�,����b�d��q$�t���[.�P3�;k�"oE�����r�	[W��O��3�/#Tzq\���*�.�o��n��FE`U�t�0^X�O�6f�U�K!�e9���g,�9G�.�*�0�ڽ��o�~�~�������p��0G�e�-�l���SJ�$�]f�o.m���o7y<�Y2]���P������G�xx�:��Y�>q@�����5?[�Y&�1��a"�H�"z���}�'(���0 �Z��bhL4��=�-&����9�5�mNL�j D�0��.I�����K2�߉�f<6�iSF��Ɔ��?��w�[�_͛��gx����u��(�p�e�%���Ĵ�E�Ng֡{�}�7ҕ�#&}�{Hr�4�٦�FOeh!2�p�q4��L��3.h����8(��PM 8h���o���q�&���R���X����l0N�2��x�F�u�h@5�U|Wu��:oX�:� E�w�YLȱ���Y�@��RBe^m��qO�&�&��ކ�A�o���t���&Җ�5��-��2d?��� 
�� .��0]#\��f��s�*�s�Z�J��f�%���+w�1R�pǼ���E�m���x�jK�wZ��������Ҁ�W} �]�:A�H�/��ݩ�	R��c�s�4�2���	�J�֜d�o�& �a��n�vAmO��{j~r�E+���L>��Z��g駋��lۺ���p�I�����>�MCI[�>��޺m2S&��.-N���ĭ��aIXlUj�����g8��н�=�/����r0��e�䢰���e�WɵF�}�ׂ��&��ڸ�
��]4
�a~+O&��F;�X�}���.Wc&�͌	:c:�%��y?ɍHΓ�s"2�� �U�0�p2Z�|O��gHD׶���/�&sA�_X@�����<	��}�,ͣ��z�U(�T�qBo�67���� ��q��W�ŏgZR��ך��U$T�B��@3q�`fz�U��Q����a������D��_B��B��!�T&��1�s���-<M�`�;�l\+��l5��u����r@?1�e��I[E��8Gh�x��c5er�	W!�����w��PV(Էg;]>�fj��-ǒǤ�� c+|�Tk]z��~���m!�:�#�??���_,��Vʏ���k��?�`Wo)&�8����!�|?�y�sC^�{g����4��UrxjvX��q�\NqNRd��RAq?w$�"�5��x��@��ϕ�4�wyz@�E=I�v@�Iy���6��iX(uQ*Os���?���I(�ON8�||��b[� _C���L���&���9F��-�4p�bl�'����?�(�Ng)/��`cf&^e�˘�P�o(*h,ʀ��j��v�K�x��<�l�\�M�����p�>"V�Ʃj�~�i+����۫c�%��p��yI8 �22��a#E����8��`M��k��D��_��d�V&>y�����m��-��pL�l��i�atd�W��g�����y�����&���b��2����f)��-�e-&����a���o���*���7l!!�G�r:Ҵ���S��*���1L�ْV���Ns�����~ҧt��^yAh�B!�?W'8ۅ���e^*�ob2�@�[њ�u�G���
���_�	5o��Ed"�SZf�u��l
��0c��{����O� ��:G��0�?�����1�&S��g�����̭ɻ�c�V��%���k>� �Z�]DU,�:�Mʷ�b�.C�&������P�oI�����xz�
O��ݱi�"4�$�=xm����-�Z`n@>�ю������G��O�������d�j�<p���4j,S�����o!!���l���Q]�b Wo�Dw�>���m6��p�~i�R��&j]W�@��*xZ#'�aŨ;�*)F�y0��K��vR�)hr8��L L��S@�b�.����e�u5S���A�˖�	Q@��t���fޣ.�3"F� ���������&?;�8��,2�
B���,_�˔��v��E%06K\��E �Z��c%8����4�(�h������֧w�x	���|=��)X��ĶP�uS���[��)��ݜxfC���χ�B_5��O�ED1m����t�`�B����o4e��bu�������k�ԍ'1>r�i�B�.���ܿ��)�MG��/mV�>`2��8�¬�,���_�{{m�KS\����a��X�W�5A�Z��8V�Ń
G�d�Ct��������)+Z��� `[GG�h�kG}K�s�E���O#��'7;���`I<�r��;�X99Y�*�3���~��}��Z��͎����y� �ğdW��<]Ku�����"]��Fn �;+�����=R���߃W��v�r��y�rD$��iB5�'0�Q�p��ʙu�~�K�!�Y���w�Nz�M�4�eya8����z�D���c�Qюm�)�Lv�Z��f�B�kv�`?�"�ڂ��C�%�Z��Tlw��3	��Jî�b�w<��Mq	�����E���6�7����ݞ���xѥ��.QU�,��Z��7L�YG,ނ4lg�t6vr��
��%�g*
+m픆8��_q�<Llh\;�)�h�lMa���q�����ng��RƬgX9�!���=�y�U9�7;'������1�"�!-W�B��]9B�F����,<V�4D����$�x��6�F.��] @��^ӯ���IB��]5t���7�u0�*�<O�v��� y�Zr&��cy|?��_��A�h7�cro6��4���'d%v0���2ڀ��z~���G|�9d,�~|aK`�����g�w�E�V�����'L�F@��K��)y�E ��������  ��·9�/� �_�>j�=(%+��Q�S�A!�x���(����a�/$��ﱼ��d0͹x1K��x�E��Ch��Wi:��u	��I|1�����mP��U�h�p����4�;��C�$A�z�_?J������Rk<ݝ�>Vr�<�Pn����o����F�ٶ�ȵ5��{;po ����`����D�N�c����K�?�8F�\~Z�뽞8m��J�8䳵JI����k%��B���L�D�F�<X�+���������Zr�l'�+���_���v��J V�� �;��p�']W�����{��?/�"���X�6��ol�H��Y�]$0����<��-�G5D���^��=��N�},{���x�b֤��RSړC�mysp*�`c ���'�|�i�g��"U����K�wZ~�	��)ZD���F�b|o�xCW9�=A�Ez5�5%\�^;1<�/��˸�{���H"Q\'�,���}Ӽ�k�f�n}�8d2���9Su|�u��9���٠7@>V15�� {D�ud.���An�Z��/_^��!*Rf����6��Q �7��dV3_Z��o+���2� �E�L�nX5�
F���$GE������zZ����q���@ �`�0�҃5L��5Q[7n�qC�hZe��J9]�
��V������Ԡ��D�#�7��%�rR�E04�YK���מy}�G:�/�m��ziC��)�4ڥZ?��f��V�L��CK$9�~QJG��?��Њ#��K��
1�=��B��B�A���_N�.���� ���L���6E��P?U���T��C�&?�q������vHq�~<1/Rw��$�T\en9:�SZ�<��&l�a���]�H�����SA�R��*M���m�gF�Kl �0��X!�����o�����d���7�K�����\������/��s8������8\���CvL�9�	�SuEm0�Q-b� zwG���V���d\N��n�Lw��H����W�K~S���ϣ568]q�Wj��Ѽ�,T[)V�{#�FG� �^Ұ�6�FP|�u⬿�iuQ#����K����靡����uG�$�eV����U(��uS!�v�s�1���Ey�t�3A�PR������V�R�m�#�?�-�����A��j�:��J�W9Vu��pW�\�L�V��W����:��D�������c&~ۡ�`�:�<y�eK�P3+��ב���$���q�o �L!�|�>�2�WDU<�Rs5�D27⛐�g���|������QM�>���Y��<V0�.>���0
D��R�=LL��f��h��x�&�E��S[��NJ�͠!�K0waI��z��o��Ǚ~E'�[|�"��i�N�QC��i3Ș�ZO�^�Oڹ/o�fOl9n��e��G�ݢ`�
��t���eE�4WA�
�EW$ߡ����JL ?v�b��[]�b �����<B�o���~X�؃G�\���F��L�.��GӢ3bѥX�F~�%F�����p����GK�e��[�8��%��ƾ����Շ<g��N��K1��!�+c˜ �8F�5V�����P.����3��ÇNA�����mi(�6d8�h�^τ�Lx�_2u��Ĵ:���8}0� �������3mby�����Q��â����ɫm��*ܰxq�C����a��A��3����}̽ϼ�h�[ts_����6g�z�!��q��A)A�Wq[3?��Qn ��>��Ô`"�)�C�F�,�+��Q��P��4j ��jM�`s� -��>���h��h�Jy�8|7^M�"|���bY*����n�*��/R�p�f��$��(���מ�,D�ςcX(���4k�L��b`^�UF����MӶ�O���]�Js#��e}�7�W2 ��TY����n���q'����4d��L�E@v(]`ZTl'9��,�F�&�Ф�T�xͲ��-��l%�wS�)ē�8i�f��pkS�����|�[2���>X��b�!�]�g�ܓEWx�5�|ӑj�4N��HY%�V@�>xB/��z�r�'���b0��𪊞�܃u͕p1R����8����îe.;|���������+��
Ѣ�;c��'T�Ig����b�6;���fn8��!v�wY�)t�J�ƕ��%(��U�)&��R�땚P���q�s̉�o]{��K+��WʹS�xJ|o��،�;�2u�]��G�9�U�nJ��hD8�����4q=�p��~&�P�S~���cwLc)�@ف<t�s��T�^h��ǚ�fB_�$I	���=�;y8Ԫ�k�^�/��	!�pC�枵P�=g��l���l�t>8���X|�������S�l�̳�&���S�z���@6;+hSMo2 �#�@"�q��Z���W�:��H}Q7���zg��+*��Z�~
�n,aF�=�ä9����P��0�}D6T�0���1 �{���ˀ�q�[4��lR5��w�y��t�/3����6��g�4��SQ^��;
4l	��W���{���-�2�tPʇډ@��N���^Q�4�촰	!u�V/mi�@����X���c]��0�x�aF֧�)�q�w����û������l����C���G�C.�h���/������$Q`:�}�DAQ�h�ʟ*-���(i���X�9��#���H�	�j�!�ޞ��ɢ��B���Ǟ��j�������K�*@�#R;�*�G͈#]��� Z�#�.@;=����N<���I��=����m���
g�l�TW!1Ye�a�@v�df;�w�U*��L��"$�O��V��!�ɯ_��K��Wl!�*!�4��C�@�3���%'�kl����zG�0�ZC1�E)�ʢ��-ӗ'CY��݄��J �����#�]��d_s��Q��g�J��g�M���0��5ٮ�r���b��V�I��$x��������݆�� ��=�S��G��l1\��3�d%f*�*_�B��$��q ����3ާ��j���%�UM�S�~�I��|Cy9�g����yA�s����C�X��JM7��k���
��)�"<p�� �����Z�N���BCAĐe�^̙F���Wb#�Xy����MoRqu�����9�l��{�Opo��c�G��[��p�*w�/x	�bY�w��f��6�X�]u�������u���9��B��.�.��տ�_�mq�<�߇�/��PQ��!w:ԝAɔ����+1���d`Q���B1�{fOU���GsG����4w�	�E5�{��dq�v�[N�I�*BW���|�rc��x	��b�ҪQ6�?NE��9O���f���:A3�ƞ���Kk�@y.��,�r �����d,W���|)��X����˃J1�n�n�iC��*E0��B6J��]��9n~���x�,��fl�L�z�J���u�7�8<�ˁ�PU�kz�#:S7:����s�!V�]8���-�Jӭf�A�Hj����B��c�ѹG�,�#��!
�7��u��81���غ5�T��sL�9{��3B�r�6���亩�:]��{�q1b֝<\%�Ia�D���d��m��u_/C�˴�3ۘ�LM�3(gh�Jq~�2��֥yd��Q\��k�K
��'"�7�[�U7�Fd\��v�U�ɌJQ)�Lua����[Z�@�dô��+�6.�bc|�<;^]g��!��x����%����"��T������X	��"��&忷��J�C����,���E&H�.�x9�]������^�r��s!�#�{��=�L��U�/n�b��EpM1�s�V<;;��0
��f��"23�c=I�z�2�j1D �!�=�*��76(�ǉk��SN�?R����_4�px ��T�dl�H���I��C�Oli(��eK�hQ���~7���{��Iyƒ����WV(r����ՠo�3Q4b$8����m�1�9J��?H!^�S��#Aj�wCSG���L����7f��~�A@����%�
y*��/�⎥P�~�S��F�[@FW`��|Q�3�XD�!Trm��"'��xO���8Lټ��Ph��
��Y4�D9p�	�1�8�~ ������ut��U��)�1�؉�A5Z���Z�8��\/�Lo���aT�)�c��k��g��9�kOx�
��3�5�C�
���ƺVKe��2	sH����?�0���gC!f��ں��W�k��ǡ��8����E�'��Ev�0D��[���&-���p� ��K�x9[ɚ�����i컉t#�a�&i,G@�P�u�	]xo�3�3��ʯq�F�Z�ȿ��*�<�'$\�l���Q�U�y�Ic�ff"n����u�+�+���)��f�6�ZA�&�9ƀ�f�O��@(��f�P���U��U�_T�xX?j	��ϬReWw�Mf⅛�}Je/wb �W.�c끌��������]Q���/Wo^(��S'��BqO͢�|��C�FyK�E�#�Q����E]�u�ĉ,��@�[�,HNp��Ŭ�J�7DK�$~&�;6�9B.�P��ma�%F|��ܒ���i]I>)�N���{���ȱ�)C�9�c/JRt}�s-[��F��Ռ<rH�n���{�����S��\m�B�x� a�Τ/�V�gW�Z�:�o]Vu�1�Б�lЙ�����'!�б�7ڌS�1܃��u [���O?4����F�N%Uy���JW��cn���b���4%���62��������츍H���6�z]�4'�Z�|c�5��G���FR�]���`q�C$��̠=gI�lR4��q�$�;�f�`�	�v"s�A֩廟��I�s��2��X/#��ҟ�T@d�hR[�����2{�H�r����y�:�!�<���9��~�� ���<�3��@(ԾZ����ݒ]d�n'����6y�E�U�T������z��M#}^A���+0��F�o�_Qvj�r�Tm%�1 v�c~	�5K
հ7C!�_���#Ule2Y�I����C�	��$}C���]������ǀ'`����r����
�j:�q4�H��+i;s����+����$�S�C���
��Al��C�L��{�~��^T ��x�da���,��F�A��P4뎖ƻ��m�T�%|p��a(��z`�d��_���x�� ��J}�q��(�?s�>IR�3�0[�wfs�S�`�������J \�D%S*`���`r����OαI���?��<�l��|`�i�
?�٠y��MP6b�%�����<�*h�"M �Z�3I��+_�/{2������,��s�O�M�;A~5��)'M9Y3�⅞ ��9��#j�����g$/Av#0���(>"A������Q.���. �i5���eËS� \b~|�x2��*T�Vߝ�7B�p:}<�A��U��e����tOJbG��t���~��4�r�D萒11!��[r�}o��uSX�Fn���J5JE�?B�g�c������u�ڈ�0��0'��!PP��rU�PP/�	�Z
�w�)��j��Wd!�\ۧi�b��`aL�8_p�*B�O�|Ǡ�0+m�O޴�6\9~wj�H|�He9�x�P��ϣ_{��( � �"
��'7�´�0"Z�Z6�˹R����1�D�1,����o��
���!z��~�:�e��*��ni:Ia��	���b��dh��%JwM�6�9�s�ds/z�͆v�@*Ub;���R�tπ�[�㍢g�,vY�%���F�_�@�%�X>��'a'��}�-�|����~wY+;�0��RN���f��L�;s���wY��~���5�@�fh'��O�C����+�"q��b�I;�t,J4�i�R�������+>lۄ���NcΡ����EQ
|���P�CK���}u��b4��FD��n����>�Z���E���E�)n;�"����,��$��x��QB�xa3�Z�
a�3�8��wT���M�����t��1�ZK8k0���C4� �b�[p��ޢ��^�:�e66��b%�y3y�0����,�#Q�;^�������U��̢x�wٿ�]ٝM1c��*y������
?�/��OԔ-.�g�,��>w`��m�@�tM��G��z��D2��d�uɏ��kq*����]C|��]/YH;�j��ٴe��BE}�;���#'��+��^)�Q/;�ˇ�X�a���3m�(
H�S{�=�\����,A�~��DL��R�� �ץ�u����yV�L�V��&_�U\����ַ�F3�@q��j��ͭ}��|�*7C��o��o�y�$�b�}�B^{b,O8�)��4�*Q.�8,�Ϸ.��]��$��z���E{�AP��ʧ�(k���H�,
����̩rtm��$2}�� �Y�2*.lE0[� {˺$[8���_��c�>���S3nE1␞/,�O�h�1ޘ��r�Q6WO!�N��E-�oTΌ^���C#򲘼�]�@!�s�.���6�u�3n�R{f#��B����{��b�\3�JɻN>^$\?|ʤ���%3���`�JM08+4�E���[uL(1��P;�W˱�g���ҿ�C֧V7Jc\�VɊ|�z���8�A�DY�<���wϠ�Jc%�X7ϷQ�F��Pr�7�m�KQ��!���$9=
5da�<��j3�Rg5	csp������G+�N1���5VĞy��Oz�h)DƎҖ�y0�U	";���f���� �@mܙ�\8�$ud˴�D�0�<�ÿC�7����
k��5��n��ӥ�C�&� ����[���Q�aP
x�çU�=���s ,�]�����v)ݨ�oĚ�8!��V���T�v��4Jgg+0��6���H�߃�o4�p��"Pǽ(ׂFDd�ƻH����b�	�� ^79_RO��P$c���$�X�u����+NV�a����������꠩�x<�,�xJ����r���q�Ѓ�����^��ө�C����������ws�Sc�i���,�R�h���%�^QPjN��U+�Gy�a2��J���P&3%��Xw�"�qAi��{0}

��;bK3I�N�\jD����-�&W0�x-F|%4A��B���4L����G���k�
A�|��< t�1��F���Q�!/��]�d D��1W�xjdS#Xq�<&��B8��
|���{9M�ȡ��_^?Ap������Ty6�aҖ)f�M��j���N�7�M)g��ֽ*������g�Ս�M5l(��p������l�aaep ��p,���C�M#�腪���=�7)�GR ���*���e�eLg�yGd��|}6�d !$��Â���@���zޅw��D����^$V+���9��E�Puy�Ya^���w�g�i���]��\cbmP ��)�*�a�o(�9�!��b�x������t̒������De'�]Y��1��9LxyU��p�>s�5+�3x��j��YD<F�#�ߤ�p��T;b�F�!;���4�<\���s����kԾ��)ki���j7������b�HN��Z�Z��ъ�0��ݕ�����0�ҧ��}�Xn�ۢ4�[@E�\8��_7[�|�!3�qi~Q�EJeS+�ٿp�.�����?S��bAIR;��SE��۴ N4[��nz*(�G~��7g'�7(;�\]��k8x�Ï��9��)4�����U�T�a���e�|{,��#R4 E^��2PK�V��Jw|�������. �/�P�=����O`Gj�w��F}J��/n�a��6cj�%�dFx���F�Y�7d�������G�/&�3�Bn��H���ͽG��j����^�=�OK>�>~ݮrC�B���� b핋�Ey��
v�#��X8�����cP��/���<��_h���܍��N��Պp�� ��@��m=h�ߵ�n?o��R9��W=�����������TU�*� �8xO~���V�@� oѵm9�G�x��4�6%d$,��)�&�MF��2P�tȻ�ok��I{u���K�֊�6W�	Ӕ���p���מH��jlo��k��jN?bsô�5�'稽��j�޴B(�~�⳯`��s��Q�H��"H��
����&N���u�!���V��G�~9m3~`Gay��f7�]�Oq���� �}73kXE�-��)�L�0D��s���Ԭݭnқ�f�V#���J��^Tn�%%B%��g-X�m��g�*�X��̱�|[&u^H��T#t�.�Ϋ��T0,tf���7E�aK�h���a��y+�ȴ?��7"�y�+�T{Sx��@�IsM&� ��0��h��QC�j���ъL��8�� ��MȖ�b���#R�:�w���|��[�|�������,�Q���Ҋ��bz����ї��p������[W���U£z��Ų,�|+���6��7q�^+������ޱB����;K����sa�E2��<U�@@�h�r7��N�ֹM���W�ɣnS(V~ڰ˰x��3�Rk���=�q�@C�{��r��%�ː��q�$s�n�F�0����tbo��e�	(��?l9��W��=�O��r�u�I������Pr�]��x�b�)S�\��!!��w����YN�H[��#�ր��M�`13A�*���?� ���LVE� aZ�l�+tFl�\��n�s`�~���5��
�?f
é��z�����a'�Tb��0��}��ds�p,�3�Bةc#����4/�%�@�v���� l4�d�hA��?�3��u>��i���VK	�`"��	sE�6��kGH�{����>�e�H,`�`@�)z�^"��Z�����Θ�k�!�ā�d�L��jt�Lq�M:Y(襧/~`�	-�x�R�l��y���I�c�UL��]d�9�����RhiB$s��6��̿��]�!�����A)��<�!�qP���*g�����)`����[4��"1�k�����{9�W"�qSeA��bA�DAZ����jy� |���ՙ&A�օ�i+�7>��F1�}�f"�rPvi�0��Ƀa[Z�#\s�āXn���B`5��?4��9�wv�QCRf����2���i4�L�q�迆Maٓإ��
����}g{(m��w;Y�T�>$F ��|��.e�`��eC]�G��9��c�� M����\���h��( <FGw���C�Acq55��^�c�n[�Q<k:Z�cD��ʘr���J�^X��jzz���^�K}�;��
8, ���� �UZ:��o@�$���G&)�R�6�?��>þ�u�q���\t�2�I3�گ&c�-]�o�d-Y$��6��c�7�KD^��2d@���lkgl�M� ݕu�����Y�0�'����������I�Zb��CEq#�<x�u~G��[���)� �N%'t�#�
��u�d-����E�tJ�(!ӃB�cj4ǁov�LF����0���R��*յI���Pw��&��j*>����\?����q#h�����#v�pдH:��3b}�����s���m�v�e.�X<U��	6a�#`�������?�R ��x- 9^yO��o;�H���y)~cR�J8�eᦍ]G�[4b�]�����38"~]��5B�h�<��� �1Q�C���g�8�}*�`{���x�N��o����H�UmD8���$+>.�	��(�;Ɛ5WN ��]uj���h�G=���횑���>�6o��}]��Xt���S��;�'#�`���H��V7w����p��i�Y�tO3p�τ{�<���z1�T��~��b�/�TK:)<�6V���7?�T.�BG��&�"G7!�*���>L�2wG�5PU,5^PM�](��7H���=E~�n&�퐷��%���K��E���9��w��߶�s��/{Ȉh�&ۂ2m�i������S��f�fF;z9��9����J�f��D@B���~(G%���c&3;Ϋco�	Y����n)B/O���a��*���/9<���.�H�r�]� ��������>B����P�#���Vu���eГ\�"`K�6��O}&V��6�h���b��k��0���`�T��u��h�	��zݯ5����B+H�!�#pU[��\��Q�T_X�C��h�+����%�V~|����/O?��>"��ؒ�$��8%���	?l�|�9c[��w���g>��>�����C~�������\{>x�ѯ=@.��oP�^�/��[���wo����?u#�`,rֈ�#��L����V����J�������W��/U�Nю������|��r�b�|�t��G�����o��L��9�av8!��mf���n	^�;�ƈ��{D�b�!5HlϏ�o.$Q;y���խ�"�9�����C�+�9�3H��Tc�؅�����6J�4!q���q��Xe�a������?�ʱBx�{a�k����K��	���b�+�|Y�b���?R�����-: K���s��߼-��W#R��̝���u�e�LڏYUUR NOsms\`�E@��bSɅ�#�B���Yhw��������Ӭ:�ʽ'Jmd�!q����Z�.e'�GO�D�=��*��P�n��S�(�Ɏ�b�z�U ��L����0b�q���0?�+��Z��Pb���u���F"�k��z&�4��IE�{�=̈́5��Rן/�G��{���JJ2��M�+}g��^��t���KOV�pfFe���WJ��P���+�2$ԯ.��ǜ=$K�P�r�� �[��MR	F�G�?��O
n���T���t�;o�`S'�c��ۍ*�LA{y��&&��	���|�6M�5�lo���yWʠ���P�σe�IS�� N�]��
��~��O���c��=�Ҳ��_ �BU��11��! ��JL)`�k�
�߾h��r{Pr�C�i�q����M+b(r�XN_9�3�.e�'{�./Hn�A,���3a���]߈g`�P���;����h�[x���J'���@
����?�km��U����+U��G�!�yUc����F�oj��ٗ�+�l�س����U��!	��D�&�BV�s����æ��׭�b�`A����s�l"���ЈRV�W��kU�o��K�ð&�sֲ��l\�d�XQD锻v�����T)�����LȽR
*���ݷH��7���ũቶ�v�U�`rV!���a̺��EN�,���D��0-y��[~�^��đjB`q�|wz��ٖ��$ԇ��1�@�9%%:?�>��Wt5<�s������j��"�����4^�wJӆ.�	�V 1����o�G�E�nɅ�D=[�*L�۾#-���h��6�p�Ɖ�Aq����t@\�,*������,<Gϲv�q	|�z���,H�NK	�M$�
�����4�\�K�k���6���*i��嘦D�7��BTI�%'����9`.�U������=p����gsZ�F�ha�]��ݵ�T�H�C�]r�zެ��z�@�&��3yV�mH��k&��!4�J��e�,_U�p9�ժ̬��M���Z0c���ې��F��X[�R������)�[�C0�3�dRpf�����b�#�w��@�Q�
�7��9��=-�$;��W�˔VQd���;�!�7������m^&t��k�27�?��G�n�Ύg�b��	�%����j���z�/NG]6y�3�h~[�{ms��3G��ͮ�-nc�<ϘB_	\͟Z����xK׽���M��І�}�^-[
�����7��D�^
�O�{��� }Y(�hͿ��.p��}lk ,�V�E��J���t	j��>�IV¿M�����Ih��3�x:�9�����=I�B��q�e_��:����֬p��@RUc:��v�j�;���������F˛憷��^��
ó�qu%nO
�OO�xtu>dX�5Z�|äd��w�{����7�&�1��^u���@-4��@�Q���|J���L'��&Q
��?U<��ד�k�g`x���O���J쵝"�����렊�w�k*���D�TU���ݐ �_~�ԙ(�ߚU�(�n�Ad�G5.�b�;�Q�yjBmm�ŵ��%L_CB�-z��o�h1A_/:&>�RG�a���{-"��psh�L"����ݤ�
6߯j��C%�@ƀ��¥ ��O�n����s�e%ʪ<�. �c�ܭtzM�Z�s�O�Q��?^�x �A^}��o���Xwы���8��Y�-'���:c��X�^R=�y��h�$EW�)�x��q���=_:�Ӝę���,u	�N:�$�=�ab ���l��A�s�� ��P�V�u0o���_�|0��U8M"�@���]��uv�X?�{@�
l�kg�
���n,3<3l���ΐ��l��	�>�8jy��E���ul����Z�?J���~�~t��%���=?���nn$�-�_��f�s�2��rpd���F�I��ب��ƏH�I�-~��JƤ�<���@e8r�ͽK���,��[Ӝ��ͭ�P�������Eۘ��bl�\̀��q�i��Ɖ�ۋı�V�J�"'��$>bqG����hw
a�to@r�{�*��8�9t�\�Y�BTD;�_�}������A�mU�~�!Y������\��K~х�g"����X�G��35�����Waj���uξ��>��?HE��)�/;#a�ψ(h�$��	^��Q}��ښ�ϊ����L<[��ۮf�l���������ε�n�I2	+0��y���'��i ��q;V�M0@H\�C�D���H�L��v�wRK�W�m%��C�Kl����;���j�،��~��g{!���<	Y�%��6$��A*)H%�E�%���4��>^���r����R�_��82�b�V�I��,�z�҆X�����|P /��r�oU��^%����z뇱��̀T��g$M-m����RIş�.H䋇B�F��j�%��Ca���I�ٜS�hH��hHZw��g�f����u���7�1c�*)��l�А�kR�|�P䴽����rkv}�;f-�U�'���)��έ��>Ȁ��L�g7&�Rȹ�,����0�9�s���BjS8�h!�Vl#��eq�]�ѭ9˒�Ń�J�?����(φ�My��Hح���?�ڳ^�0��c�"��t��V1�!���TK�i5ĆyDx��R����������s�uKK���=��J��� �ɸ�/d��?x�׹ ���,�6
t������䰡�*�-h4�2w��qS�j7�;�mh9�4z�h%d��ԯ6!�(�K��W[�����1>,(���nV�?s�xh�ݰG'�Á�g�U��CR*HjZ�m�u����m�֪�b����8f.�LX�_��"�L��-^֚l|� ��C&Rbg��^n��=��YB&̃�x��ቮǭ�9d�No�ש�a���U	w;g��=��ڀb��a���Sg�h[x8���W��\ r�Z�Y�i���.=�"u����,�Χ�\��_%]��F{���e��||� �S����0rB]�z�t$Y��>3-zE�r9�_C�L��=�h�cQ5@7����_�O���V��ɍ�^6{�ҿ-`�p��5PY�����O����~�����٨/��oq�>���eO��w`����s>T=��'e^��%���߭�㯈ӝ�tU���p�M*)���%	s"7�Q���k�A�:M���w�o��3�6�B}$��(s2&/���?ZeZ@��kJݴMS��Q0�e	�T
K.�v��
ьKN}Eٞό�^�a��]��!/�v�!�������?�)%bU<�'6���Be�]E��B���/�Ϋr�j�DN��ո|e���*�����V�?��o�8��D��y��w�
o){&`+�ID� r���Z��o��\�凬�o�fQ�u*��5�������f|~}
�(/X��IG�O��Xc-ߠg�1�iYK�Ƨ���M�	-?�T8��};F0�tH
S�(�8p�5���ԸM����G�6 ����gA2v��|��"���.`�G�`�h��ۙ�Cv�)ј$&�% �[����5H���`���g�l��>(���zc4����ŉ�dj�Ûm~<yڥ�ka����rG��8���߆W8wh�Q�x�A[>A@2nM}ۦ�Rt\8Q\�'Ap��q��gNQ�􀜈�p|\[�:D�W>@#|�R�b�rZH�o�ܸ ��cB�u�D�a꾧{��>-�
���2�b�F&���-�*������h�:=9�W|g�gGa��`۹��!Y:�%Uӆ��$!y�D&;N��zhɕ����l)�з���}+C;';���놲z�]���s ����d��_���M%#��\\v]�ZT��m�$q����/�>O��:��F�P^@��y�|s6�S���@¿�s2���$v�>���/��8��pd�R��C��ս�W�	p��L�3�m�f۲K`�xH�RJ\V·��}7p�s|���=��p��� �Q�-�*�e�jB�5����뱓)�����cY�rsa��*i��e n��$��*jqv��9xd��=Ȉ�B�H��b�,�3��X��o0� � *���9z�\-|������'8����6��L|��c<�
']Hf�>�'~ڃ��ɩ��%�16��Ȱ�K&���C�������rDe�$e�Hu9��:�����91a�Ae��t�V�C�m 7�졳����b�r�\b�j+�B���
�:�3M�V�a0����o����(X�B-������N��h�|Zg��"�~MX̼o�$9ǡ�Ke?j��V�Y��dw�A��Y�Ys� ��%�S.x��m�j&R4��� �p�?=��������U�z��gDm���hK�<[�Q��,W�V��ޙA2���A,,�A�sA��UO�Nzi�W3�Ψ��������t��|�S�<N�볯�\c���'�Y̺�1<�!<���q���ۗ��M���RE�%c�4����d�xa��I"CW�4%��1�s��6ȷ2ܜo��Gʲ���1��\��W����Bآ)��ؼ/mrbC+��E��j��A�(vuim�~w���C����O����ط	���R�Uq7H�� �W�~��nˢ���$Z�+x�K�]�?z��`z��~��e��x.e�֋j*����9E��ݦr�H�cp�L+�#���g�?��l;��tX/ZCG$��#T���k���	�E}����6{c`}K��G��A�ۼm1�P\�;�9!�E*X��@/���V	qZB����ʇs�m�.����N�ѱ��o�P~"N-��!N��0x�[���s����zr�DD�Շ[������bnq�ߧd#�x 5{I���L;X���|h�j���H�qm��]��F����$�,k�I6�����ŗ��\Y����Y� Ɨ/����֊�X}NWh]׎�o��w�������<!5�O��^�-���<�|�9��&נ��Pʦ��oR�����gp�%��i���&�l�V�p�Φ���Mq�(���^�7�i��hJ���J�����ʅ�U�Wz__?r�*����w�kA�������zƸ'�[�'�m�E8�n�,�h��ƧÍ4�ܡ�=-a��ߌ���F���6�'xIr__5Z�EmԈ=��+�LW������<���uK2��I�j��#����:����z�oX,^f�W�@�n�\��d��K�	���>w@L����ڝi��F�p]^(�:3z`c�S�0]1��E��@�����8�9 ��q�F}�E���ٕd_$��9�(s� 3�4�F�Y���r�-ZR6��4�<�{�M܅I#���Ȇ�i��Yi��W�]��yng8M.��������Pq�2W��-=�x��
�m}� �C�*³����N=�l���(a�����Şc�%��zKU�m� )�+�7�<Q��\��Rl�<�l$#c�X�-{>����yE��)�>
����8��.G���f�e�:+��e
a�fx�����B�c�<��J`�
٥�ϋ�������G/���U���<�q�wl�yd^���2P���Bt�L�����:݌H�*�Y�7v�X�L�!�@�-��SG� ��GE��;�|������<)�T�C����R'OXA /�	y�������(�k��&��_Md�d�P�#w�����o��o+�nJ��=��H�u��=�7E�}��,�x7}�4�Ӂz.w��e7J��+����]�(�
���v�\	�'�F���͠��%�};=ч"��w�!K��:�x��>\	���\����r�r�e���R '׷�WH����#�l+G���� ~�����6yk�����.�'/�$�^�|�,��LGn%�J���Z��h��KF�L̒�}Nΐ��j��: ����Q�x�R3|�7�/�{�dUS��p�Z�qs:L�J�^�s!��5<�"�{%ej�u�M�M5{��Fd�	%q?�o� p��S��W@(G���P��G�R3S���9�,��h��yt��R��>��T�b ��U�-�cdp.�Iz���a%�2"��௝��657���8R�UM�����i�@���f������dvDM�Sc=;�|���y�S��f���6�޸>�����z��b�g}^�y��H��6����7�뮗�9�Y����3c�
��9��0����/�W���j�:��V��7��H`C	��R�
��܋�ԂQ�"1/!���Io��H\G8��?)��.�
��jy��-B�c����
,������H_zQ�`Zu�_�iX��y؃D�KS�2ª���eϕ��@�Q���IxZ���&s�[���jl�T�X��{�n���=�E��5�ˮ�#X�'ăx������?0�],�����F�_�1ڟ���8�jGC�p��װ`�cc	vV�4���is]��B^�r������1�l�oG��L���Z����Y�ۨ�mG��l��#W(:95a�������*�`�H^~g��ĆU+}v�3x ����uAO�䅓�:�)�J��^�w�8�~8�p���E
��'ʫ&�Oj���ø�Ż*�)f�a��8����(���$�7w �@3Rֳ�1@�`��uD�J���L����������j!3�k>m����r�����p%�"��2�}q��";;g��'w���
r��|����� �I�6VY���_�5�k3����L!j)�Ϗ~�Ặ���D�4�~��������c��5��Ly2�����+1�E���Wq�s	ms�.��$���F��8Piρ�����T:v�+ġ�IUIJ54M�`���Z��1)����`; U��P�v)�d�b�w8 ���_�{��7�~B+l��sQXF�q�ñ�$�,u�� ~�J֐�M���>O���M����XO��Ye�u�E}8�0�S�vncz]�|	Ic�Q�sA��g��� �]�{A!�_�/ � ِ٥M���ӂv�-D��|F(�fn��#�5d	�������Χ)�!M��'c�]��{Qd6\��sLk�0m�j�6
�y���⧳�jpȑ�;��o�k��Gf*�&��h�p�+�����m������SU� �_�g�E����gjQ-����uF��������(��fl(k1�.i�r����?,TE> ybW#�>�.|�g3s�����/�����c����Ec�=�Mt�,��D�n��U�p�f�0^S�i9��/ؔ�n�C"m��w��a�U�Ek,�4�Zr�_z�]�q�L���Qd:�z AG��Ǯ���I�^,B?*��V6�5p���m@��Ң7�#V'{�=V!�XF�#z������������S�S��鷀�ќn���*�QbU��b�DY4Cx&�Y���
e}tF!�8pM�te(*`u\��~��}3>��1��2���DW�D�K=S}���)��m({�<��PCvW;���!gf$�b!���R��'G�Nstu��&�������ښ�������I=��r���g�aɵ��A��`y�Z�����>��Q���l��E�AH�LT���{�Fu�~=L{�ǤF������f���F%�q��C,�"�0�|�=����Q.��ϭl��¨�t���S���-̀�-cFZɄ�)���«�i��V��I^h{䏀�rM�<�CmG��a�v�Z0���-�G$������e�%h2.F���~=p,@5��㋿iJ"��W����M8�6�]��J.h,��U��[Ĺ�f�!d�0����N@7P~��a)��;�p����w��5�i�����U�J�� r�u�#h��e�&��W��6.�݃�!��(�Ṵ҄�4�}t��H��a,3J����^=��CX\Er=��y(-�:Ͽl����#5���2`����;�o�"��T)�WTB=6�"�%�߶9�v/��!y�=1�gW�O ��
HV�6`��Xa`9d��'�Z#>
���.	��)2a� +�p�+Vʡ|Z�L6ht�`3��0_�U�|���GQ�8�5 �A�D�q&2fj����P�L�b�U����qհ��x:a�3`�B�ԇZs�2�/*��:^�;���݀�{;6ɸI'�5p�H���~,���-���:���ÙFUÑKՙ���p���RFØ�>d����ɺߕ��2u����w��0�^_]�� 0���&,I��}�IXy+��rJ}�zt�*u���2�j��W��N��p,�\�HE��g��^.<���FY'b"F��
�����0�u��aJ2�=��2��t�U�˚�ՙ9�;q$o!��&&cr��Ji�&g�.���2N��[7v�Gi�=��K��>�����-{������4<���W�A���V�0�"�R%���sV-�I�e|4����K�ֲ+��}��$ �`�8���xz������y�����?O�ko��!� �**�*��o���$7]��P�l�!�#8�����k�ʰw�������]��.��@P�Nj�Ve��3Hn��+(�i0�^���a���Ycv i�Xb��p^ܒ�V��C�e�F��Uwp�j�hg���?�U���x?��G��ɯK�X�:�Ri����Ă�����Z�apx:�FӊvO:./�ۭ�aF;�Wq�[��yޖ]>L��=bZn��Bb����ܣ)�����4��i��$��R��:�k������Ň~i1SP��g�b��<���,�҃,��ຎ�틊э x�� ��vU�b�C���~�$�4�Dj��W��[���0l�p̀���K34����fΪ2���F�+�	������?]�!Է��zu���<""�%`I�t�zFf@�.�7�T��}����p��+����6�H0�BƠt�:x����gg%ދ��BH�ά{�,�r�~3n~���V�7��9Er�03�LV߬R1�E��|�[I,q��yG���b��=�+a~=o��ڽ �@�q��v�F�/�	�fk�R�h�(�f�� }R�������U�U�V�T�R=F��	?���R|忏bL�?|=�����<�l%�?}�B^ ��Sd��WEA���[m�ĪO��ޣ��'���%��n�'|p�1�\��ZY�{ٛ-y��j�r~Sbx����=����y���Ŕռ~�x/���3-��H��Г������r׏~˙N�D�͵}�ĳ��-$�d�J�0�V�����_r;f� @�����
H��7I�u�r�7z�*:O7<K񩲈�ymj08A=ls|�!;�ÒuF!"��3���&ig�w�X:���{���;��L������Gr���ﱀ�^#�kbB��,��N�Ͱ|��.qg��ld�pt��.���ھ�D���iVϦ)��wP��RB��J�@�9�	�hDLǶƦ�!m(��;�v`'fp��m�~�:���	\�W��������..�1���0g�����,�k�-Qz��2���1��|�1k5=�,i����!��0KQ1.�p���dز*���+x��>%��y����s�Q�������hq͊2����Rh�<-.ZC�G�? }��#�`ue���G���(��7�>�\)�;��03"�s���h�>���y�5����Ҹi����=�f��C��S%X�ܦ8�E(}$m;��v.���÷�Z�T�IcE��O�ʁ3������m�Yg_���M���C#3s>߄R{����!�?�n�q��>��*�r+G�X��,����@�x\gh��� f��{Ϣ�	�ФI~��!�%d��R���,E���&�����>ߺ��t#�1APE�Df>V�%�BW�4�{bf��ZƂ���C����7����~\ď7�U�K�J�y�50[�J��]������V}MČ��
d�UM���Z�H�f3�k��k�5��
�S�D��B6r��[&�j���:��tG �,%��P�;_����ZI�%�5T>L�����<gE�fN�X��3�F�]�,G�V���Q7Pe��|@�Z��-ے2����YHf'���~�����INz�\O��."��9�T�����^/���1p�"��6-�f�ɂG�����5+����+��Í���o4��-yT��_��	"�{~���H��}����"�IK�������r��-�L��X.S�mh0M�!�X�*w��<(�`F;���N(�O�</��):W!8$�a���'�����u����5����mZ���(/��-�V�79�L=L.K� y��0q���M�iV��K[M�,e%1���$XC�{��ȴ_c�%�#xBG�|[�%������}���x�NV-�t����+�� ��"�?\n�G�f`5XFI+x��3 ���^��K%xu�e�]��Ĭ6�G�p��Oه�Uc�1���&��]�&9�߫�����ԙڽ-�NZ���[��!r���%�X�.���.T�u1MM]�Yy�>w�1�L�QS$���(�yz�XY��n!�a���3OXp'���l��M������'`�[�v�0��0���	a�36H��Z.�&u�_|p~�zRL�����ܹ8���	I}e�L#Wao��9�������Q^�����{D���5 U����У�Ґwy�.E��V,�^��༇I(��Y1��ZY�m�ȏ X�B�m��d�w3��8��}Si�Ƅ����ߐ>� h�@g�P�>�S��^�|赘J������C %}���P�h�31���T-od#:u�8KT�*�J\:�vI_kt"E�����R8�_�_-�\�Tx���H�0���%1�;�yH#Y��Ѝ-����{�ڜK^���(�<��1x�Ջ�.0�A�C J,́n����Phtq21ث���~������M��>n���L!x%W�cpR��U��zy�1��ܝ���An �9�=�pԜ㱻�@|vs�
������ڇ��A-�t����+p�Xd=��Z���z]Kc@A���l�4/<t{�6(�}�}�H�.bo�9殪[�RM����-d�)d�xs����@8�N���u���K�^����������ޕ����֕�ˮy:�xkU/�T��UOH�-��#���:��ԼidS�z�[.%�6Kɓ眜G�j�/��K%q�v�7(����I�ٸ���no���a�95��
�a ؚV��{�m��J{�����
pۺ���N�8S��M������%`���/mr��<�E쭜E�`@ʛ*���!؜���	$��k���6"Hk�O��8�W��y/���=���.��]���r�V\����:)a�Òt� �t�ۦѲ=-@2�^Q�S:��������w<Z��IɌ�c-�����*�[�b;6%�4�B�l^������e�1v�F�Z��|_����Rt+I�`��fU� B��O���HAL�S��{Tҳ`�\77q�Y�Q�4����	����@/��d�P2^��)g��s=/l;y�A��%����iI�70pK����:��ꇍ�q7�QAB�Z��+�<*��7�}I��vق\�ә�b�Ξ�eZ��[���0� 2;�k�Fɴ�e�,/����Hc�n����nZ��O���Q޳|^� �ʙ%Ʉ�U΃�f�]Ac����)�,��c���i�s���|���)�4��I�Pԙ��}�{��[v)������8�����%Ox��N4�� ����e@�N����v[p �[b�s�Œ���յ����Rƺ�iM'��2Q#'k�0V\Y�C՟{��ƒ�(_众��UR�0I�!��s��C��tn!/�W�yL�]B_��"���9�׬�>�D���C�eմ�^�`|a�=��M$�4�W�X2���5(?ߧI��P�S��iFH8ƸE룲B��AgA�ʧ$�����*�[z=�BH�emr��O- ��8���R/��_����i���r��z�<���Pr/�o���i���r�»�P�&����J���$��̓�D��0���/A�n��<n'��(��h���k�eXi3,��s� UK��X�E���	HH�M�b|^Z�v�/���
��Ah`Rv�_������������:ۨ�&�8;�a�3��#���N�C��ek��{!��@H�bqNQ� h�Kakg����`-mh�+�G�Ɓ��x��^��5�;�6�37x TmY�|t�ŻM�Z�ꢻ��S�\H""+q���F�x�f쭪�gpd-Ϫ�&�0��\x]�^,B�
��#���|��m����ND&�F�S�<�"�X񁌣��z':rEBg��� ����k�$��8�P`����j��z��=Cm�,<l�1���A��n��׮��sX�S`B�I�����s��&[�n�"1���&K��M�� ~�hv��Ƭ�j�(6�.�J+]��C͠������X�6��g�傋\���76;�>S�篤��f]�q�h���b�8S�F.X�d݇#B���8ۨ�?��pxJ�T։"=8��F!�l�hA�g�c���Q'?��횦N�;Fh��.�X�!��7{��b}����Z,�\�I%�ǎ�_ڄ�/w2�1�}5��,�.S|��W?)�E1ƌ�N0�?�-�hi��r�� .)�|�.W��W��������j�`�n� �k�u<4�Ye*-5��Z�|F�v�!@��!Ƕ��.-�cB{�����tQ�_���X�j��Dk:�O(��|N�L$r�J���%��C��e�'��Z>�� ?(���w��/
c6���,�ȝ�v��)Pӛ��	�S�	�J0��nǰL���3�;����<�����\c���eݽ�{��&�* �|��!���X�>�Tɹ�m�"5��6���&�$�D�eR�4L4��(*+'U��r��ݡ#'Ɔ��[AU9�w�AHg?�@���<�+�U�@!���i�ĺ��4�q3�'�D?D#�jw����J�=3��s/�	E_|���Fxa۫�N'�6��>]n�ko�p�7�uz�X���YO{3� o���9�(u�W���]������H/�o@Fhr��xavZy��ܨ�h���0}g �$PH4�1��M�Jv�B�q�;�j�_Ã��"��p��$��⬍�co�~��Q���~�c<�! ���{a�ze�,|�ha�0?]����ʅ����M#M�e�̥�4�
w��u�_ϟ�Aî�hB ޔ/1N�������I;�%S�H"k���i-/�������p��光��=�v��$l�_�%2����)��*��,�(_0����>Ђ���-y�S��}-;���a��F^�ް�_���������ߥ�Yë"|H*T��F�/�-"��4ypq'\o��f�q��Ǘ�|� �nBN�~c�<J���o���d��N���{I�U�?�]����3+"{��v$�����E�A���y7]Ӝ��x%�6�kl�i�X^2bGf��WV�'!�ھ�M�+�e���h#�h ȣ/�Miy�?P����y ���2�E��tu�=i^���q�U5�t�� �R�pD���G5}�
�Ka�+��M7'd���!��/NI��0L��V`��J�I�k��p����T�)f.�!~V�W��^�O�uۂ�� ���͋�ޠ$���p'�7Դ�*�J��{��߲Zq#8vd74CN	Y40��#��UC�Θ-��Zt-/q*lgj��WY}�嶛U2� ��ʦ�O-o�����,����� Y4��N��@����7�Z&_�b4߉O��'�
Ͱ�[�+��4��v�)�d���kiF��`G���e� �������N_�d�@�9u�\C��fr�[r��Ұ5��\BdvZ��L����E(���F�2��GZ:(�Nժ]0_`����T�la!ą����� lS:���!��pk�i��kq(���R�/�"`]�}3���ai6��Pc���G֩��`��Y��>�)��d���Tn��ьf��ߋf����XJ���3
h2.�#�5ȫ�1N�Z6�_ 5�p�H��%�e���--ߑ�*wsX�Q��X�4�)L� �����cM�C��N��b_��C�h'�3�.<���A�>���ZD��^P�����l��K�y-��6.��z��e^lT�~T`W0���h�Ga��v9��=I�x���e�c��� e�|��W����/�'ж�	I��mt~��+mfD1띱F��1��R�ml����P�Z�f,xXYD���?-踢��H����R����=��'�Z%@H)�*X,�U=�$���ݧ��=���=a�I!P-�"V �*���0���9���mв��r����W0;���z���d&
�75k�R+s�Sh�}���^ ?|C�d��(�b%d�[�\��j�D���{UV�xc�����cmG�0�N-�p�l���#o����9�R�r��-��������Y�U!>-A���z8Pt���ʰƔ��KOYG�$�I
��[9��3�LD�X��Tnӓ}*�sS!��N��l����A�+�o�~��JV8���x4~�[�|�bV��E��������K�5��Lhp$���JCX����˦�L@��Dā3�@�&W���i�K\�aD7��6��gq���D��U�E�|�·��-gj90>j���M�wEZdA47*�[F�Qa����OF�Eǻ$��\�<��@�����)��,	��\��e�嫉y}��� ^X=�zM���{�Q3���?"_�[&����c�@��z��l{`1QC�O����t£24� #Ūy�ki6MՍ�'"��dx����Z��t��J�]qS�|�m
�+�t�{ى����@��I���N&��S��xUd ��j�~U��L�6Gx��忐��Jv�/�+M@�<R��Z����z$��X�~�'����<�Gw�������i��%hN�i���H���>���4f��l\���I�{8ৄ˦���]����!��m~]y�Eo�>�_�8Y\X�m,����,�J�-7�qw_K��웩���ü e� ��o������_X�⫅}[^I9p�������}5�[tK�	�%Z�������Lw��NL%s�����&�x�����,��w�t{:õ�j�g|�<@d�s�rv`Ӵ�&��K	k1[���9R���GzO��2�?�'N���s����)��=0�@�K���7� �X��ѐ63�:�Uqv���y���2���/�e`Cy?j(�x}	>��Uү���_;�ࠡ	?�e���+��BIZe�n�d�w��뙇 p ���Tk��-{!Vit�>�B5¼�5K��f|�h6/%��
�w���s�C���нy!���������c8�����(����������Q���v�H�w���XYf�X�����^��&����#E�E���7���TZSP*� w>����z����'q�E�9����sH����i�{�����HO)��={�/�y�	�ݐ��UH���1���g4	NL/<��Vr	w�&y_�b6�ȋs4�ص��Ziٌ)|6"��J z��T�23�`�h#?�h~��~ �y�I���{���u`2)����a��"�ؔPGn��#(jg^�[D����_D |}�gt��.%����gI�)�Rz�J���O*�&�V�����f�L�yN����}�#v���;�t�%ZY�e�nU�l~Y���t%d�/S�|��7.f�I����ƙ&KLP@=�:�������Z��������5r�T�{�y�_?�	N��t��4�h�\#ڨb�{��FL��TȅD?��v>�ث8NE�J��a��o�\��� �-5���+�Xӡ�����;�B|�'����+*ܟ��_,7���S��y<_�9�I���L�@��D4v���^'�'��w��1ՆV1ik��K0��x�Y�s�L2�����r\��?�"��}}V)|'�tA䪼�U�K��r\���,��.fI8��ߟ���d0���:�i��V,t@�����Wn�h��6�g��,��7
��t��S'g6fV�:s������h7=��3ݵ[�������|J�:U�Xi� �,�i��h��I���&vd���|����&��+��ɚ��DQ]�W�����
�\vuy<��'���3y}/P�lv�?�ۓ���$W~��5���ޯ�Z�Mb*�G��!��Y��9#R�	�~�/����B���x�_-l�J[74�3�2�s���h�ڝf�?�ƖDTB�ږ�L+e�O#&e
y?"n3I�_���D��
R�1���Uhh���M[���dM��� ̀M��9����tD:��f�dzT �������x)��'�w��ˊb��ڂ�U3Cz!����J�	jg�͈��1~S�x	`�G"e�E�P����~fΒ�������t!�K��o��͊Ɠ�7�J�"��C�Ȩ�������A`��U�\�{�
>�iќ��K?���hc�z��_+xg���Q��M9�&�QQ�M�ky}�	Ta�)SӖ���m���+����/Vg��Qa�9��L����W���QR�4�搤�:~��y������k��r�;b��cx����?G���s1���r�V��l�KD0��)G��� B'�l����>8�����(���k�S��/���$����ε+yÎPXv%�ʿ��!�Lm[��㟞��m͊;�����|��1����������
Q6Ƀ�,��GJ�笎V^+В�<�1�^�Ϝ.=��)��I�_�Js��cQ�('&U�)�v@��F�l�i�	=��Ē��IS1��4�K��;�,�{�G:/G�G���[祿����Z�<N���O��b��R�X�����]��W:��a�P>��ʟӢ�I���3.��J�?8X�I�7������KC>ZN��Z��炢8l���Ș ���i�qז���M��r)��ۏf�d-3��y?��)�LP��(�d�NH���i���ged{���n��4Ю�-�SX�G��4�a� +1(�X�� 
�`X��lvs6�fmm��ڒ���Ö�%ѥQUL�E�CȔH�+m�J҄G���[%_���N�H��Q�=���*by��I�	����D,ᆛ(F�qz���(r�&A1�KMw?��� �!��#"�c���5��y�ոl��t���K9�A]a[�������LYh6h:��|�s�I��l����d�lV+�G�6tH�d0���!ɖ 0�]<0V�M6S�\ln���T�V��lo�w��{$����I�f����B(��'���כ���%j�)?���&dĨN�����Ĩ�2݀]ip�fV.l�X�$��Y�7s��z�ǃ��	\�h�Twu��3��>`�Z�O�PN�s��L;���eHˠ�P��e3rw`��ԍkD|"�$p�e�Dp�8a`1+�w��i�D�$����Tފ��%M�N&�"g�����k�ނ�2��FR�۟#AR8�E`w����ԈTk�%��vrS��*9Zs�]���ʲz�L&��#1�Czx��c�b��Z�4)P`��F�̔.��ݮ��+���c�~�� & 6=���S����	�JUЧͅ���r�׮��&�L�ؐs_����AW��\[G���ya��pѥ 7�Gy�m[&��)��za94!J`�Wf���֫�QN��~f�l]�?�XD_�C@	ZB�ϧe��7b�6�_�b�W�/�䴒xU���_�	�]���e,V4u���KL�.T�%L�����7n�4�����k;��]��d��:��?�Z��qe���5np��[Qv�I�ƥp
v~觓�n�n�m�eX'l���\�x�� _���  -��Bx3덽�e�A�7�q�ɅO�)�����ju�q�.��c�e���zwb����U�ĸk<�̆4�8�<��H#��ݖ�D���gPc�;��2b)S���G��j_CI�>z�K����v���9����6fU.|�[Req�3��(�!�45�u�Ӣc/��_jc#Ƕ�-���2���P��>RA8hE ؉�Ai4
_w��h�t��4�C8�+@���
�~o��uO�>�C��C��=7y�@#�5�RÏ
����5�$KF��G�0��M�Q�(z;w����=N����`@m�MB�Byࣃ��$�O��|Ӌ��ѷ��Q��_5��
��DT����S�[�O�q�v��8��j�v:X5��+���@t}�O=�[���ˡH��"��`�EMX) X豀&_��W�AO\�9�����/����i)񡁬��o_�0�]=D��}�|���KQ3�X��7�PՎ��8���rɊ�?� v|����#5p�����8���@P������Je%���y��z�h��f\d�J�	�k>�IV2I\��b�S��x��#$1���Hv�-졭ml��5���'��7�� �i?�-#�~mn�#y#��F3kER���Z`^�n�r��{����%ui�I�ړ>��/Ef&���G����gg_���U��3�N���/��DU_�m͕D�a�aPz�л��OthU�v�����wҡ����zK.��ɔ����]r�L2g���CQ7븗$���p���v�%��$t���jDbLɧ�7l��"րķB�w
^MbOQ�Vq<�{Q��ֺ�z�o������f���KI���쏅;�'@cK��Y�_}�i�!{1w��k�A�N�7�̭��@P��XDR����Ɯ�k����	F
�u��d����\��8xRF����Py�9_r�����qaZH+4��*>�Ml>.�f��x�i�0~]�I����>0��M��:��>s[`W���߻C���Ķ<2�hT^8��=���f3)��@#�u���j�)�v�b\/��h�3�c	w���'��>���'�<�T k%ٱ`K���ޏO"�T�tDʹF"3F�4َ'�Pvش����7��x�]5���E(�	%\��P ˂����lS1�[���z�w��a�,J@�U9����ǅ}I8�E�ۿ��$4�̡���Կ'bŔخ����.�V֒����Ky�ՍxQ��W��n�|9�C�y�u^��V�)|<�4m��\%Ƀ
[P���ҴQ������|��T�i<�=���t�R-�)Q� \ڍ��q�җ:r��]�^����7��T���%��+[�u����3{��xL&~!��8Å<�O�K=/H�5 ���Q���;�i)2�%���!a9��O��3��x[ڊ�}6�C��78�Zy�,î|~���..-�P����,�y���^$�6��Zw*;&2r 
&'�X�����t��%nI.>5k�I�a��v��,����q{��@��&�7�J�SdN�`�d��_�D�C��7��P]��}����bL���va�#�Zu�d��E���aǼω�tU�A3ޘ1s���^w�>&�p��������O�ݖ�o��L����e��&�沸kKP�;�ҶYW��j`�bB��+>p�-._65.6��%��:[�����j&����c�8*et{��vW�G#��+qX;�~rz6�FO�6[\I��Y*�t����֛~z���2K��'8�d�d,�`��s���UB��l����k����>_J)�=�Θ��ګ��Ա�l��W���0k�u�o�P���c�vN�-��0�(P�e6Y��pl��x6�͆ڞO9p:�(rj��H������T�@=Q	K���7G���Eޚl(E)_�5�ܖ���hҢX�N}Ch����jWjX�u�(u����eǌ��Ǜ"�����F
"�Z�lZ=��x���$a��y�	^3��unu�j��3��;�T�p��!sd�̮-�T���l+zF�~qGQ'�y;1q�F��s��ILƈ��km���,�o��7e�SΗuI���
4-+a��n��昴����l�u��7�h҃��08t)3O���-�p�9����Ѝ��3$����J���e�Є����V�`l@J�i��iS��t����#7>q-��lP��iҨ����	��iج�t���ܼ�kݯU2�'^} \Ή�(J{�^z$�R5�q��xf�HsL����Ĉ��H.�]��������c��]�������%���88��U���z ���ʞO�M�hE���h��=7r?��\�C�a;[H�O�l����P���`��O�y4��!XS��������:�JTZ(�j:U
"
����l-�"�3��֜����9�}`��w
�;���j�U�?��VDw�VDަ���d�Q���%��~�9Aa���x��f�H�|~S������"~}p"_�4bT��3�2�G���q���*x;���.�km$�
��.ⴀ5����"g�z�L����
	�j�^�vjk�}&��]�=���;+Kk'�+��q>�V����T�{'2,�E2�f�������0		���C�r�E��%5�7%Cx��-8Y�� ⢫e��9Rk!�i��/�Zx4���@�؀����fA�h��_��	�ϙ=&�M]j�W��k�<`r�fC�(�-Xk�NQ��;��C�<e�~��/�ҝ��y()�,j����eќ�Ap�gD	��G���gg?�A!�s{���&{����@Z�x; 04���Bm�v��}2+�Һ�6��2���J����;�h���ɉGe���I����q})O���-�v�o`=c�]'wT�\:�T��p�DIGD����~Oo~m.��Z��7񽺬�������I|�tn=�7E�t�sP�}�&�����̥��a3fPsT��:�CRe��2U����m��A�r&d;��@��P���Kj ��1�L�IX�\�O�*�/�U�[��,���}ax��H���q/��d�C+��k!�H��U1/��6ǔ��:Gn+Y�\���u3l�ω��*	�sM}��*�[�ȝ�S��%1P�*pד�G�TD����"�f3ў���gH*-)-]T��B���`e��W��+��SfSAߘ��MǫW����Ma��*�n�L��n�����	�=�jъ���jhʍ��]de1ԆeN��5�ܦ8k����5�s|���՟	{ s�O��k�0%���C|B�[�q��U��ʆ�A�m���PU�PB�-����wE���9��n�q!KC����\��j�tB�\�:vV�O�^(D�@��1�|�\�ҝpl��LEwL7uǁ��g�w'쩈��~�B:?�����H`ש7�%VPv)δ�.��G˖�M����Oo���rH���z��(�q�G�ٕR4�5�4��	�t�>�
T���-+��'-5��M>}�1��� �م��uE��Y�s쿹���.|W����}3���I� #	l	�.�b�e0�4�o&ŧso�$��D��0�M�rX�M<Bv��$��>~���bRi��K ��K5 �'�[���,7���8������
�7�$�<��W>��)]��^D�1Y�k"`{}����2g�NjnQO�!�%`�"be�tݮ/[�W{�B�!�� ����tp��9We]�M�t�etX���p<K��+eR���ñ�)W�����>Đ[�2��#
i��J,ot$����M�{��N�m��ׂ��&&��)!�6/�ȕ�x���[�t��?h�"!H��'�
��������k��gB:󯢻P���J�x(p���?�o����g�uO�v�x�ݓ�l@ު�5�����)=+�vV���O Ot��͵4�$�9'!b0,R�A����q�.=�>K�&��ߜ���v�*_���?Ӹa��0dP����)��o�3��f��ś����yq����b�9[�U�BSI|b?��<G��� z�uzĀ�M{4)^���47��	�Cl���_�I	��'-�AB�0�R(�Ê�"�4�DCG3,�E&��Z�&�|]�SZ�r9���e��u	mV�a9J���πdd�]�<�oY��^�/K�ăؗ����lL�"CK���AW�4��:�ᚁ&��p9޲ϭe��q�_�[E{�,CxhϚ�@/y�`��V��?�g����@t����9��8�:�~y�ښZ������W��������\�/��V զ��
MT�CȈan���4�J���D�DF�_N&[fl���c�����.M�Gش��mZ�m�i����B����D�C��߻�4e�wJBVfg�4��Ș_}��N/hڲ�OiT�喼T�b�=���l�޵,��� ׎Eya����.AQ��)�Tns�E��i���2}utLmDɤ���{I��wQ@��x�CT�ؒ�������y����^~��I#��RR��YQ涧�_���y�C�^O�8�M
ZO�	,t,�������2�Q~}W��bŲ���b�.Mo���CF�gK���u�]˛Cwn��lW���X�:o�U9��ܕgL@������ŝY��ocb �;0�.͟{�]U]���q�����5��K���
|U`��D�!U奇�'���&ڤx&@�3.�\/��`�̏4�O���S�$bE�3�6���z3w	�K����,ָ#c&�י�S��%�^A�xi3�Et��#93���,*�w�L+�M~��6��8l5�7H�q��2�xO��jg[�7�#7�F��J�2w������K��l��?N�Tc!l�y�!�F-����GV�UO���;�&L�"�d�ਨ�m� �ρE]W�����𸔭[&\]4p��OaTďXE������膨�f����j���CH)K���N������d��Љ�q��L��Ȓ������	�D��M��24�4؊
�WQ/d�M
��H���N.�����e�`<�e�����%x�����oT�v���{��V���#2t���OѢ��3JC�� �;�39%�O0��z�n���`����*_��sX�g��|�>����s����Y�
�;��t~X�����XK�pj]ڙ��r�6�u[�@L3�x���k��]�} �UX��M���S{�V�{��\�Jo��&�&��'�z펾�2-���3i�<g1e}(Zލ�O��*��4캣������H6/��To�`z���ۥh����~7��ކ]��hZ�ftL��N|`��Lwh��i��G���k�ٜ�< � m���@C�qԭH�/,a�F@L�K2��Ξ䉥�vc����Q�kCZ���j���{*|����(���4���z $7*6j=����zR��i���zpX���L���AsBvR�Y��e�jW���E��)�'C�2�'䡶��k�:���#LW�G�m}ٞ$��yd����<�( T���
��.<�*���9�j���WP��b�$�t`�'r ��UL�G
��OTS�+|?f���;����s�>� O�|`��$�� ����6�C's�qBʫ��^;  �VГ���mj:z�r�ו;�. q�����?�'+
��1	��<"^H���A�a����+V����w6�;G)E3���ӂ*|��>?�����~'P�}�C�<�;N?3��a�ݜ��Q��A��T0U�N�����m��r�x(�x�oq��s�G!�9���[ �ny�#Cs�!�ŏ��c��a�,���>/�;T��%������4�w�3Y�_Gꫂ(�u�5Ҫ����>^��&i������d'����d�앥�#�}����xpn� �5��FR�P*z��xn����<M$�3w�욢Emq4O���b"�)��q���YWYQW��W��n�@���l��#�eq��Xh��V������U�v��d�脠12fH�i�[w�y/ʁ�g&om�vP	4	~g�,Ŀ�[�8큃���B��������&Q�̝R8���ယ
�x�4�E�D��4�]�����m'�o³�]���{׊��'���M!� l�+��>��6WsJ���W��k�BTtڢ�����`�nr�}��'����V�� g̚��4�)/`<L����4������$��yc�d[��u-}�1C-�?׈��9�S��i<�x{:�0]��KLqn�3�R(B�K7P�qv�C3�+�m��L��^}3�G�O�,K#�� ��)�}h���iS8|>�ʹWRG���L\qjQ�Fe�D�gz�lc�ӂ������x~x��l�&��.�������}�}����Y(��@$Gah5�+�|5�Nw����l��'LI�#͋+�dnR9<A<LK��[�8����{E�E�IG��5�1cPZ���d?-��a	N�/������'[)����jM� ���v����(�S��;��Z��?�f�|~���KќUW}�	`�F-�h?yM��ʮ�6�ı��E2��,�.lj�d���&�׶�K�RLf��L����KE��q�G���=�s"��۲OE��e[V/K�/���!�\��$���q��k��{�~Nv�`݁ٞ��J��[�� pX����a�d2'p�{	�>LnK�/h�7�br�tUt{͹��wc�NL{�hJ��f�;�Q�aH�c9���!���c�W��5N����e_��®L�&HB���)�V�3�M�hɧ}%{+�fD|���"@+Օ��H~�Gaa�#�4[�#�E�Ɏd�ܶHΚ�1bjl�35_}B�5L�2� ��� �,e�l�KX�!����[��jCjd��u,�&��q�\�,p�W� �s�.�q0�3(u�٭�`C�^TVf����g���0a�ʪ�7�<⻄^���~>{٩G]~�dP����C���B�t��k���ߤ�%�z�J��3��y/���/r�6N5f���D�ݢ&-9�p~���#Y+��Gw<	׍�d��F�`g̶��h�����ٽif��й�Z;[�"=��o)�����@|�x�Tj���)����T�,�W8�Ij��vؐ"��B�%�i�HdAgIQ��N���^�x�/w����?�	��<��~nzh�	���k�Y�h��U#�=��d��a(��U���	x,8��U7�P�y�-��R��o%����@�]dU>�35pĺ��҆������".��e�SS�<��9�P�5[
sdNÃ��J�,�>W��li���۸�/��Lف���,�e6)�&�ߋ��P�*3fX�9\�ɿ5�z3�u��У�1���{�c���<�H2��юH��AH�em��)�����9��EY��4v�Q�i�p�$^��U@��gؿ�wׁ�Z0�H�	׺ W����l�M%�L�Wa�M�`d(iK
�0̥�[,��$�R�@Wr�I����q��^���<�T7(ڴ���-�9�3d*�߈ː����>��>�3;A�����<�9�V&$�挻�y�㊎��?غ��j0�e�Y�<�T`�<q�4�.��T��s�[`�_�n�#�FX��XS|�^���0�v(��F
���{m�w��|�#o�f�y�vX'Ŧ�%ou>Ѯ�)�{,Y6�ZGʋ+�7�̑��n�;}@j��~�B}򤾪�]�c"�{��
dT ���咎��W��.��#�0��shCS�с���/�ܭT���P�sL���Dy�,��36�� �6e���tk̇_�]�&5�q��q��}Im�]#R�����C��!Ws��FFFexS۰y���o:{��B��G�}���z;pKV��s��Etx��O�`��J���VW-��]b=����u*b�����b�+w�j�yy��'m=�ֶċ���Z�LM��b���[�9�kTc��/S�m?-�\en�	d!����g����C瓪F����?�3G��v�:g�+�vѯ? ����e�ƙ�6Vc��(AeU�C�<O
��-)��n�Y�_�ù@�$j����{�ژ�~��R$  �9�fs��[���c ^��.-�Dx[��?nUPM����^��Cdc7ݸT]������Yy�*�����C�ޝ�X_�!\yŖ��BB�>����E�
R�7yуRj폄+�?�ē5�Sp������1.�oT�"?��>
�B�� /�f�����,��8ɂ1�xQ��^^ju��8��A��#6t�]�D��tʒ�7�V��	��w�`� ]wF�q���#�%�:} �����8�,oO��슳� 9�� �8��c�+
�KB_���2Ɣ��;�c���)�a���sfx��W���]UE*����&�.v˛5{-����k��׋� 9(#*"���x�X��U|Q���3�I��4ٝ;BSB��si�8���eY����
�Z�o��b\p$��řlM��D΀�:
Q\Y�XmM=4�JI*|�}G ����`i�:�g�8���T). ���6>x�#tXč��fU<��v������Kr#�6TI�� �
=LB'QU4d��d��yíaE6�e;ǻ�G����!x����Iّ�O�B�_�=*#a/z'�TG2f�RȌج�����X�����7e�
��̩>�B�����-�WT֡L�����!9?��c2�i���ػ�������%T�^�~��^�^X	_�3�M�� '��Q(=��K���\F�v��C�R#O���g����W��e~Z�C��&�ڕ|֫Q���	�A��0�c���H��~$q�\�d�r�k�����M�=�jNw1z%T�~�F�W���;М̐��䷙�v������r�Z�wz�Tzjok#va����jIhY����P�a�g�;�f��L��6���T��|�0P�I�37B֣0c����?#:n�7�h�!��ӥ1����d�"��-��g�CF��$�	�!@�������F[��%��f�p�">P�i�Jq�zp0��"����]U��������J\��FK��S4�Y���w�.^}�����I'$��� ����$��u⹴�U_�l~��
��p5]"��P�;"�Q ���Z��7���ͭ=���b���骭Łn��L	� �pn���1(q�=�ۖ�λ��f
��.?��K�i�K��Po�\�{#�����o�S2���98�>	�����:W�{4|��}�Dd)�y�짩�� F�[�_ ��~#k*y.(����r7�����1������l$ME��R+�b�r&�*&+Yq2���cO������> [LyV�\�'�=��ɣ\�hT��*�����/�2�o,�j���D�Z.���b�>�����?�Ρ�(n�G�-_�L"9� �t+3�ܤ��+�o����3�\|�?�0��Ai�F�m���}4�K���$h��5#9�S��*�_���^���m(���r�2\/]ut<p���j��AB���r����d����__��QF��<�R@+hv&,r�����y ����ژf���C�"�+��������ޓ'v���59Vt�U�6�Mu���P�[��ſ�^dˉ�d�~��ǹ�=ͣ-��^��^9h��V���%A~o�ǃ_t�`�K٪V�tE��[��k�V�(g;}`�*GF��Em�7>NR�,=z�_�+�����MR���\ŀ�c��og�*�ع�$�G��B�2���X�zm�����;�w0$_;�/4?�ԡ��?�s�>Ŏ���#ގ��������9����Q�U���J��D_��I�ӯ��\�p�0�s�
zW���%熾�7r)��*�C*�0������0� ,G)V�m��&��e�-_�۬�K�[�>e3��m5EsC��ԯ�E�@�e#)#����єD�@%�RM��ӻ��Т��;�XX��"���~{q��MS�Ʌkn����m��hZ�^I������RkCnׄK���r$���������_
��)P������P�ʎI�M�e-l?��w��Վ�0�_�w��ZY���oM/���,;^Ɩ�.��0�"�T��z3���=1]�(9���a�m����LxM4�2�i	��l����
�ޗ��`��0�F?�.['�yI�K孖3͑;'S�`-�eu3�4��������N�Gw�!grW��l<��o����S0���o�p����"�6��n��O��Аe�d�cfN�W�����tt�0��o+��s���Y�!^�w��|�<��(�d2�B�Uy���+K a9Dg[]A9�ɪ�G�\�A���/�◊<�am#� �	兤r��F���d���έq��^M���qi��<	�]P;F�FF��R�_e��npkp�}_��%�xMQw�!�js�luJ�X���υX��U1|�����p�bѦ!�0	R���ZJQ���X�{<�'+����`uW]���y�(��N k�=�i��D�Lۮ4H7�$�4F��z�h�GŽ:R! W- R�]���M{V�����bR�*?�"b�V��)�F�^�X)\ٞF� ����L�Q��ϧv{�G8��C<��u{��C���T3ԕ"�R�� ��C	**3����9:H)
�Ѭ.���f�Dq����7�g��n�@�?dJ�չ�	�,ђ��W��N�Z��;ٓ#+In?^�T���T>��-@P噇��#1���S2G��[$�	�K
��Ro��U-pz��A�l?��"y�y�;��?{�u	D۵��2ּ�Z�ڕ���V��k@F�m-���O���$|��m�0��¡�5e�+���Eˢ���f�p��V�PcO�3@�S�ϡ� ��P;����rH#����TRbÛL͂2�Ge��Л����m���&�˹���F[A��C3^�OP�A�tb��c(¤��6܊p����	m��	V�
y9p���72I��a�G��Bo>ϒ6��%�t@��/tˬ��?�"�BEZo[��7�b�G�^���S�a���*��R�Vޠ���!f�C��'K��K3{>���B�	���4eK���҉<p�B�"
O���+��B�ף�D��e��9$�(�G}�)�+Ǡ�H��!}�1��B���t?aO���I��@�
qS�?�<N��
����6y��?�;��'�˦��I�$��R/��+�bqYȦ����.�_�_9��d�St�����Kd�i*l��-�q'��U����&0d�(�~��[8#��cl�g�M�^h�t�/`}���0P_���}���/!4�_�3���TiV��O��/������߀G��U]tj�n٢�I�LDǵK&?�)X�.��|F��m��q��w�mp/D!�ol��V�%��cq2��3�ԕJG5�h=�=�}z�ؗi-�U(ʺ^z��P�'a��?"�U�x�G)��P�J�j����Ĩ�U�{���*z������F���R�x�ɴ�~��I�s#/�t��6�̖��8vs�W�'��O97���3\�S6�l�7��m��	�n� ��V��Rw�qx���G�弬9�ͳ��i�4kS�m�u,v�6P&E�I:!�:�iZ��N.�
hw6��'��3"s�ڒ6]A)�t�놞u��W�v�$6�=�_�LKm:µw�����{LSƽ�0�4-���럳N�7`)T�9_u���=�
i�uY��� z��<��o����WǤ�K���d`}%��6G�/^��J��Qu`���T9��H��\������[4�n,+c� �!�����c!Z)5�6!���Y�_ 'U���Й�Yk�7���bq}����!1km��m*�f�j����\�l�[��H���V/R �׈�Tk�Xǈhi��3v�&�V���5����W�	Va�攲����\���Y�@�BD���e�S����)`1F�����˟��A��)�����z��4��S�a2sH�=6��a��lw��P��`S�HL��K���=41�!�5�@�|m',O�����L��͌�n���(�G��G���tN�\2�>sz�z�`��_9���U|���BWm�R��o:x�=�u�中�f�F1�c�eB�XA~��ɁI�s�A�D!���R�3\�|%tY�$���bRq��=8Co��T�׊6��z2��Zļs����q"i��������2ݺ2���]SaM�%�{I{�R���B�]�%<A�xN;�E����*��~��o�84�,l]��8�/�1ʔ
�g�s�'uyu$ ���,n�n�(����I�7�}�	�@<D8](.y�!��3�n|	����W0J߳��o���ͮD�,`3��AN��g&'�k�E��G��R�O[z��˙���,O�_��/�o�[Öp�o������
YRX��^T��U�8��5��V��4~��n�ݥ
T}����<���FYzѳ�z{�?3nͱ��6��[�>�ˑ�7�7��U������Sù7M�#���/��*��a�V`��P�3��rf���:.�A.E��}�ӏ��<	?�`��` �Qy�"�Kց6J��Av^�mi��JH>�i�X�b�A ��uI9�;t��vR����	v�(��g}�΍�H�n�gk��)H��BA1�qм��O�9�2���,�f/�����d����!�l}� �تxX��|ѬgQ�#1��������.:ߴ�:x�vh���	 ��c�w���{=9W�G�6�Lč��x��|I�2� "c+�lv�JIXn��Dy���C�C��BX&�/~�����{"62�S�zK^X-���C�/��i�j�< I���w俌I���H��B��8=�R�H���p����Z�u�+)�K��)e�ѷۂ@E���-N���r����>r�B�N�9.�>Xr�D�������9�aT�f{�i������%v�������
��,�O��i�{�9��i�-`_���vw1%��'w�'�sr[��/6�=�(Ï��ߋ���v�H2�k�g���F���׿[�=�&�����ҿ��ʝ{��!��`_K���<��\*�iO�-�_���{J�E��}�@���ש��G�f� ~&+�\1�*��ďgr��I�6 �Sz ז��_��glnd����{#�ģ�w(� X��4sE����ª��.";�����
�"��xo%Cv��S�<���H�hC��Z�_����opck�%Q]�q��)=d̫��p��N���Zi�^��ۆ �?���Q�x���5ϸ�놃l;����|%�������d>��[��zA�}&7�@�&�WE��#ghb\���b������oo��fh.���2��CG��4@�:sR聠Z S������$�֚�m<r�> �t��O��|L1������j�vR��뜞���%��'*yu�/����'��F~�+@�*��W���D~�����Zdy;�B�P@��c�Ǎ}���"7�$5.�l;GVe�������Xª�vj&�EE��R���nͱ�q�]��w-��$��mFig2�c��nX6Ea#l��~�)��^�k��u���٥�b�;�h���n���f`�Z��oVwZ��,j��z�IZ(D���o�bx��<��Y5}ڀ��ʁ�27�G	���g�	y7j�J�;P��壎1�k�	��sF�3�~c�@鍴������:�����dQ���|ȃ�d�"�����v俭�H��G;X]��s��?Z��L�:�ʃ$~�������*���_�;x�S�cDoD�́�D��.x�'�m�Z�iN��+�����1�0��)5�T�w5>�������p��=wn�u]^*��,�֪��Ա�9<�:���z,��њ�&�V��p_���e��릟��]�+�X"֨���Fx�j�N��sW���vf��G�5�(p
b�sx����7*g��/Xh/a_�������k�w�Y���q� .�Ť��X(��Q6޳��-��x0��<��(/��tG�/�WƊc���Ĳ:���:�jYW�t~L�}����B-e�^�*�FhA�D�)D� �����M�ퟮϱt!BEZ]W����g;�U��Mx@^h+:[]#���`�Eh��`ƿC�e��XL�i3W��/������添�gs��U��v���w������ЄG�?6�Hz�@�R�|��5"�@#�T�Y�q��
�@9�5ұ�3��dkr3�.�Ӽ�L������P��8j+�����F?~9���D��k=�C�q��|j���B�����j�6K6��)U.�!�ۃ�A	y��Q�s��=�ә&����b0vՋۂ�ٜ��UG=|��Z A�|/��J\�"<!����s��/��Zy�<�0<��/	ϓ�Xd��u�2�XK\pP���Q���<���N���>,K>,�`|%���|(K��,�BhD���e{I���GA�hg��;����Aѫ�Cbf�E(受2/���E?e��b����y��%��`Q�0Tݨ�;ҭ��	.za�������}�~�?߀�����@^_���R�R��=�R�H,=^b�uq��z��&��m�ɿ���7��6��, �W�
�f
P�.<����P��1�Pa*���o��A��XyI���(�����4R�?J�1k9�8��4C7 ��=vL�l�N�.!�9>8���b�������p�!~&�z�m��g�f��*�P��_����GS��:��[�<κl���K�g�	q��y�1PT��{_l����.����46v���\1�r�wR��.1N�e�wC��7��]d2��� �I�.�~<����Ȅ�+�#�8���ԍ,����G���v�ԧ��a���&�	8���G�7���	��|��qm1�A��
��8aOb�@S�����=D<�E�q�@Y��5��#͟������^@y5a&�h�Y��I~������i����ї �H|���v�Q\���%��9�V2��*1j�Q�s�e�����@��c֮���	��z;�
X���`19�����ad'{�L`_�� !{i%O�o���̚E����OS�0�^mAU �sI"v���|izK��%Ʋo��c����8^��QI�Q�� ��7�#$�!���p�-t��+K��C�1���o�0��gD���U6��~'���=pPkt��9t2}�%7�V]�w�#��Z�ȕ�⁈H�Qf��0�8�����g������@��WLG���#�|T��'WN����J:ilu^�ȓ���ʬ)1��y?gB���tFG�/�nM4z��b�^*#�!Y��@W0�d�D�pw��,��;F�t��@y�~d�/5�G?�<�V?��[J8im$ �?z�%�	bd���K�z�R���5�Z����n�+�]��b3��+Q�������Z�Bp��x6f0���gҟw(OΟ�ˮ�����DɺZ$�ue�n�(gy.#���E��t�1dC��y?-Ce&C����H\�T/���G�/R؃�E���{�T��:�#��~��gB�~���ao������cW�������9��C�E%-�g��fER�W�j�W���v��sr���𐩟''�Y4�y8�g��3����˴�;qg�JN!�-*�+K^����pIxq�� C�N!*��J����Il��)lv�OL�	lUp���y�(ȀS��Z7ros�׆9U�r9n~� [�2���h���i�G,,��w=fN ��԰ �c��Yѻ��q�#5� � O���iu�?��B)��Uy���+��:���=�h1����t�g�1� ����9u�;�z7�90|����*�+Z�q`qğ&��5�/�5�_�cx�/P�#�k�L�L��{�K���x��pɹ�$8K~�*�a�ة���K��l}�09i_s}�Ƕћ:������W\�۽�+k�{�z|b����#\f�Rc�1K�y�}W��&���,D�t����<���p�m�N��=d�Wx���>����W%����E�K��'O�@�1(*��>s^�E�Z������ڱ+�
��~r�x��W�@aFK��/
rs[�G����~7[	�b*C5�g���I��/�^��P��&%ktm�+�:E E�&Yds0�6O��5N.���f�&� ʡ���,�|�B���}.��>�[��'G�� J�Pn2�� �(簒 �86����*��>a'�2��f��n>�7���,��H�%@>��r��4vہn^�L����!�������Y�I	�.�5L�u=\\�G�z���~��dF��`�kl!֖8�d�َ_�`���@ܶr�=%=[l!�z������򖂌{31�:�~;=.�2�H��h�� ��Tؖ��5�g՛A�~։f9���,�{��_���ؽ���,�U�P��������
��p���^G����ט��ɐk�W'27!��,x9Kh�,�W)PtO~GSo߯)��ܥ1ś�@�d!ͤ�i�#�c\�-N�G�N�M�S��1����0QV�.�{x,����+�J�>��Ӥ�}L؀�C��K�Q�js̲L<�FE!���3��5ʽ�Q��t�R /��w��N��N��J.� U�f*N���l����+��ݝ���R�f�"8��}j�݁3�＝����S�7OIօ����i��!��>�W�&�aP�J0�H!+ܤ�'�R�V0>���%	f�>3�T.�u���䬕�7��f-5t���r�H�c>�xVod����p���y��{��F� ��n�!i�۱�T�����ִ��f���KHGq�<d�VB'�tb#�$��飃@=��[��Ul�}b�%¾��V�	��כ���G�wfj鼜��8��z�6�K	��9����y�X'[�%��%W�7�.�
�KR�e	����� �p		5����t+��_hQA��`YQ-�Pw���0D/�5��D��n��!6jt�]X��[�=>��/؝c��.��j���]?���X��k���
��H�sh����*JF�)�n�G�%�g��T<rX��"o�{�>�^	WS���F�E���!�>��;fÈ�VA���5��^�&�i�؄�Ǹ ����׈$���r�\�ר��7�?�8�%�-�+<�hH�����Y�dX!���i�Pk��Og���yzS��5I�q�|��>�9u�%H5(B�Ժ�h�a�,���:��.�C��N�.n��u��EgC���{s��G�*��w8�p���d�4sEs1��?��� f�cR��KA��T���E��y���
�-b�2���~l����u.���u�\=w��Q�e�>-n��[O�z?�R0v
�*�CX��Q�Ns��iq�Ѽ���i�
jbE��Nq4? ��l��Nu΁�Khَ�~u 0A�"0@g��K6�P7,�,@��zZ(��8l�n.�W�:M'YQ�}(�+1��T(p�ͽ/�2�5GwYgJ�A,���X{�D �E�Z�.e�l����h�5i9`�O��{��(�X���7�,���mL�&���W�7Y�Qvɴ�X�b�l�]��)���n-���S�� q�w�#�y�R�����e	�V�S�8�t���O�u.��k�/��{w�e����t5D	���F�i���j9c�T��}�ݦ,��G��8H�N�i��p�Ц�\�h�C���9���m���[���;4o��"�m�el�!O�S0���#ps U��&�EIW�E~��e6ۇH�Ɍ?5�m�VƳ�|�g��NE�4y�w���4\�l8BhL7�>ZS�%�D�M�}�����_��PK,<�H���{HM�"Ma�;|&]�V��G`Ax�<uy�CVJ�1�L���ַ󦴄���E�K"he��5嫂�s����Y���nf&Qy�ۭ�8���2cñ�d�	�8HB��/�T��}ѥ�Ad���#$ge�&;Z����w8*�ݔ2rz�N�u��u�|��J`�Wa�H���TI��\���6��z�۹id@!5ԡ�U����d@�˳B��<>��9S�}�p��bBi{@nl<���9�ȋ���|�ܢXS%�h�ݪ��`x<� ?D����@�;���h�͍�6F2sah��@�<z�tĭo%��4�;\[z�����D��爤��Uh�:��mt\��S@O���|�<	�̦��*	�ޯXֺ:;�����Բj�(J��h��L1��*Z�Q��i�1�*4|}KB��e����IZ����S]�����S�����ǣD��ɿ0����U\��Z�
�A\Vc?��ȵ�K����`N����鯍	^�IHE.��_��!C�S>�c�@<�M�$�!t�ֽ��$z֎^����%zɳ~�L��P<��l��Q���H�"�Z7����y;�9=o�-���p���	�z�l��|5��03)��z�=+�z��qUl�	�V�=|�y�T�d.�ү>~�R�y{�ݔ\�x�|qzU�X���1�E>��p�l�#[
a�w������	�v�� ��QWH:� #���Ϸ�Hg�vQD(>!7{F���i�0�k~��N���ZW]y��cIS\�$a� �@H4�6�N���J��L{�:��|UE���Z�<
���5'�6r�A��J�����M��I�����)�C�Li��P7�1���`l5 �#�>�&�̬Z����+z;BM~�߀�1`f�&��J����^K�{��-+����g;�߶G
��g�R�D���,�
�#��/�Y��Q�_��0�c��n��:xu	s�.�ϠKٹD+c�'�(P�*�Jb"ʷ�D�����4����;��`��`�F�H�"U4<�m��Z\Zm���Z)��S������v\rEtJ�I���UD*v{���	D���G��*t�!�?�9vԐJ�F� �,I˝0F��>Q%�&���C�X�G��]��y�q��p�%+e�OJ�dF��i��Y��kh���"����fݱ�>�m�f�C0gj���tr�׻`��|$��T�{�����+,	�"J!���ļ;E����M���1�:�mU�M�n�%5V{<2�xPJ��:0��9I�7��"�$
��H�[l��]5'�:]�����)��0�L�����Š��A��r_v3/�����I��.�Ԓ�'DW�Wo�Cn����TҞ~�%�i)��!ܓȀg��#�t�Ӟ��F3��l�/������=}#�G>��H��d�y�zZ��z�d����d�d��-��󤬌&b�p�����u������i9�,��=r
A?<�v�S}�:�6kG[�ͭQSf�uS��t�#���+��3���)<�[�'��#�x�n6���=XB�F۟�ӎ�6�CKIC�t�4(%�ʹ��/઱��q2�j������H�Z
�����J���5#�L'�{����n��/����[��܁P���E"y4\C|���������~f�� h��Ԃq����qo��܈�Er�)�d�p�$�F؀]-���Lި��{�>}�}�[�c��"RZ�4�'��{�h�>c���גJ�.����?�Pm)@�5W�k3}�Y���ws@�6{��$�B��%���V�dꓔ�?�Y ?�"7�[Oq��DH ?N'�uF��w�Y�|�$�S��5�E7�N9�ԩ��A"��6ajo,�F1V��#�L�"�9�l�hQ*�#�d����ψV?,�</�\��.g�1���]����C$����wa/J�i���d�|~2��NȇVj��r�D9a����?i��:-�ܞg�s%: %�v��qg�˫����b1��O�n�7W��� =qH�8ܛD�#��,ňFdi�Q�k=�-��.4#ur������sexޑ�%Cz�a+B�d������Vq�Ep��w]��>궇�������3� F�v�vE0K�$U�L�zhb�Q����n^Թ�x�ݙ�t>���Ok�C�d=MPйڤ����tCv��o�gq��aZ�AU��M!�g��&烋�ŵ_�*�x��l
#��䥤�yq�]O(U3�N�I��s���ȃ�9���	-���T��&F[�q������8}�r�ڮ�t�?}f^��w~���ᡰ �3�lN�fgF�����%Ot�h�C�4�%�J�<Z<ԉ@��Ȅ�<K(Nm�9��Pr	f#�2��m�Zo��B�2��B���{Pq%�[w���r'�w�� ����v��׺<nm8-��
Sx�(����Q�8�\F����s�Ŭ�s��G�ˍ��&<8�̊{��X��qǫJ$�mpj}޴u�h#It��#~�|��j��#� k�7�K�2�����R29�ī��U�[�<�wT���t��`����wӈ2��R��aQ.��N��Ҏ�Z�e�V�H���[��jQy2���%;����X�۳v��h5"#��7{RĀ����㌦�GG�:��$�q�!�^A��uh푿��t&Ҝ�E
/��DQ+��t�4׏z�d�Ω�p�=m�t�I�k�d1����R�h��{T�n³��^Y<U�*��1��@��f@
�u�\�~����A�2���H�o�r�ᬚٍ��\�k�B�H�0���I�q�lP%g�a^7�?��� }�K�BL5���ں|������ٵs|�w�n�e���)OC5=�R_2&A�.F�)eL��6z
Om�e���������T�)��^�y�8p����ݓI�y�����øр纺SH�T;\֣z	����s�J�u,t����Hl�ǿ�m��g��C���
�%=����\JXM�ͷ˵�ʯ���B�q�~7p0�}$�1����RQ����4�x��Q��Y�F ضT�R;C��V����I	��9��+�2k� ��
kV�~�\p���9�w���&�Oh��Q*SqߊՎ*����1%�+��yk�ׁ7�5��}M���f$�+��"��r�*8����B�L�\ZA󟝁��E�lV�$����|��>#�^%�IL�}P�T �8L	� �&�_"QO��F��-�z����nN����E��k���(�Ez����/�L"��N��_Db��-�3X6�_v��q��"�D�R^�5�-\6����9r����U9���	��W�\B��m��$�8U����/�K�2�9��-Uٻ�Kz�z���o���X�������ϼ�wn�t �r�	}��d Q-�:o�z+pm�x�ȕ�m�N^D�	.q��B�p
s*c��X�>G�2y)Na�ބ�r�'Ĝ
��T��݉:O��e��e(I ��0!��Յ>�Uu2 z��-���W<~G�����Қ����R�Δ����b�t ���:��"|�waݽ{kP���siEf�zw
�� �!�R��ca�o�{i)���b�(�-q�|��z�NjM�wh��J)7�, �w]�q������v�9��`�l��(�ڏl���#{V��MY쵴�mlc�v�h�@�aa}������esx4���w6��~m��)�{m�p��+���7�Nϔ���N}�Bfx�m�B��,?W��+o�"�a|t�=�}��m�]`0�|��&�X�ތl��.�{�̨3l�-��Ye��(?ю��^8��JɘT:��"`��jB|�����d����!�m����E@��j$Ig��C�q@y�j70��Z��Í����ɤUZ��H���	%�P�ܚu`�p&����$��o�ߒ�;eF�O���mM{�gr5:��O1Z�	 ���?ԃb������2���ްl��o�ǆ<�-���#.~�A����Ti�ʙ�@d�=v��
�6
~@A��.K�K�%����Vؗ�d�b��	�T���aۥ�G�V��"W  �s��pP¡��+�2΋�m�1�4��v��w���۽'@ޮ
ߢ�����l,���t��ε|�:�4��!����]���Ǎ�=8�<�>i\=��P�3I	$���	n���{DVV�J긐v�m���c��K��TFwu<�<F�g��OW���lO�����&��|j���&�}Oښ-ӻ��ce�gkѵ� <'lч�q`@	톾�اκ�Ϛ����:7�=�4��d`9j���'���_�C��ĺ�G(�^L����۵��x
]�%�p��dy��ٟ�%�f�^mARig6<����BN��BC�X� .�D���W�\^r������JÍ3�ݹ�4' {�����c��^c]��.>.�;Hq�/�g:V����G�#ݏ)n�.���oן�?X��(Lاh{�f��-�S`�D�$���Cyg ��4P7E+t`�t��\��\O9�q����K~�q�x?�4܃f���S����j��dI9��B5}���5����p��/��$��h_�}r�~�!��	ܦ�R1�j�G�C?��u�|�sꦧ�� ����&�t��0��-Vw���1���f�� ��i�,g����,�|pžCō�~"Ux5���� T�p4�[�@�Tʫ�NP��&ir*[|c�����Y�w��W�f�|V9���sZ�W▄V)��a���	U��q{�L��q�&c��Nz�.��N*ȿ�S�;DXC	� ��Ѕ��Ý��4Iq��&�?G�P�:)�iF`C�n��i?�8%�^�J�y�*���,�3��,��854nt(:Yl�F�a*�Iy��bO0��:���>���FW�6lᰑ4�3���/���`Z�W�2��}!�t����Ƹ:$M��$<�e�d&:g�H��ĿP�+g*5(Q\��I����f{�
�M�Y�a�D2D$�ɣ�Зe�h8���&����'~U���p�� c܈z��\�|�Fl�M����Q��&��k���_z}�a
1��<�W��9"�<<D�?E�)�l9z��X�4Cc�I)�ie���L�*��ŕ�TE�z3#W��\I������T+��)��Ё��	\|�!�[��o���������4(x�b�ͨc�&�1H�Xd���Sx12)�#�������N��b�DƘ	g+I����1'�&��9�8`�c͵�
�^B�Hx�1�B����i�Ά	����4k��<�2��9�'
�I\�rO�^U�������	#8
=����[���_�+�h��6��8�.f�I���p���A�����%��\�g��#���9�3�F�A�����M��=�妊�� u+�Ѵ�<.��w�K�3��D�knp�%���4LZ�]�7p�nL|ח���/�|�.���(��׊�Q�D��i^,\z=4��VR���ֆl���K΂wΛ��������N����}��w�������������7=�ا1�,�i�9FN��6h�<�����I�RT(3��><�"1������Y�E<�4"/�
��f�����Ď7���E�`�����2�	���S)݅}�Pf�m�5t���I�h2���&�g�s�йX���:�tOB�H�k�����D���K�����K���]��M���HP�M��P)B�*��_s��9/�@	9��q��nSx
��-Z�~-�}R!�Ŭ�7�8�s6��A�=�E���HCO���Q5���ɑ��q�0�>�j]�ZqH��"k5�Iwe��kJ�g�H�Θw� �����%E��I�{�j�T�&��m�q�-�1�7ӀX�"J�:v6��AP�W�|�V�3�(�VA9ߡ������՜�������:�$�tRR�³1'�]��=(��Д(<�ZL|g��}�i(�d!`�j���8�?��69�ቜ�h�Z���^����D�9G���&�?�٨/��:�}G��|�J�V��_Sq������a�A����g��9�����p6,h�M���og�ˊt��ҁ}���e�$�,j ��/� nD,XH k��l��=�^�>r������J��l/��=�srjA���mS�|��yS�a� 6þ۽Z��xp�Q���թ��d�Vx�l���_�yN�'m9���f��
zLlCC,����e�R��s&��,��q,6IP2oR `@+y�W��� ��n[�;ri�3d�"�}힦N��	`�qNR)Z�=��3Id�6tJ9���Ǩ~�#IO;�͓�R�Μ!��l�[�G���ϐcf�v�$�&�I���p�ATb�d��DFX;�9��#-Ǽ��"+�ُ��݆�d_�V�'+rU��.�����8�Q�i�}�ɐ?��jI�h��3�J6A��|�5��nE�mN9q���f�V����#��0��=n&{�p|O�`�oo��ۓ�QI��A�i�d�����;_�w���(r�D,+��y���Bbm�oo��̕��p���MJ^��
�y��b56R���|���p���PKﴮ8��&:��ӱ�g���JFN��a����+�	o4z��
%9d�p���كw�0�:) ޫ�	|���ƚؖ���tE�=���J�� �{���	mpTǜ 1�ͬ�����X�	��9���KN���k2F*Q��`]�����w��Hh���59�O�B~�8Fz�Hʟo",�e8='(r�pg�a}���5ũV�f�z���l����}!��ѭ���m������1�S^��[��#�4���@��B$�i]w3�\�R��љJ�}�&�BC�Qi�5��a2Y�X�p��T��}\ڇvja�8�J��V#��V�����S��תQ=A�bM����oZ�H�4FI���
 ��|S�z��>�%#����a���n�4�,@��5��5�<�v�"�`*Ϯb�$�$$7�"�v��!�#�Co��+�Ji�$^h���k�c�f]c1�a��!$�}��z�T,ư�B<D�Σ�߹�h�����F��+�vs�������Ԅ�ĉ����iH-���ȁ+���2 �һ����tB վ�/�%|�hGw��ô��`=�eU���z�ѽ�1��;,mo��<���jp�L�?���pTD��Vi�Sߠu�H��,q�`.�h��v;�g<ZX��}��℞.d��{����
��������-�0B7������εF>��[�,]?�A��6՚����O���5�:�DQ�#w	�?�b�U�?}���/�|�_p2pMk���l���p��
�a�,;��I�U�S�禮���6P��-~��S,��ޖߣ��� <�ӧ2�(M,iZq�&u���"�k)���`����~)~7��Y�h����	��?ǁ0�^X`���|�۸����?���آ֗Q�\��I$s��$���/h.C`[��e�vq�2l̷i��:���[�\J�^٨�4��yX�?�ړ�S̱�U�Bo�{��1v���G����mB-��(�3��F�F����}�š�F�̀�l�/E5���Q)�?q�Dϵ ����£�������"�M��	�2�������Ł6~P�b�?.~/Q{Z`ɴ�Ul���X��|�(1�ƵF+?��6xM������H��׺YY=���I�쨀�KŴ�u�+��,ޕ���l�EOv��P{�ʓ�<�L�lvZ�ق��TP`���E�(��lb��3�^��^��yk�9����"qb}n�+�	P��ja@ ֽR�j�c��7B���	�ٺ)�|�t�����.�TZᗈ��}��ǳ2�y�{�f!��a�1��Gq�6�4�Ql�s+�8���{缪@p*�u��D�r�iQ@���'<�G�7�C�xY�3�7�&��YCk��74���T1��cg΅���f�n˔u.�`�]
B��t���0��?���V�@ޡ��TG�Uu��r�D)�-C�>�Q�|��ڟ�/M��,:IN��HPr��Tf�{ٷ���J.�j�OB˙�]kj�vf�� �y�����Xro%��/׷��LκΫ�*h\���ej����!�ˤL6'���"�����cӏ�Ƴ��F�Vx�+R�K^w�T�H��#���� p���5�x�C�%ɬ]K<z ��b 6�pP"�`	M�`��.�:+�xIIGV��,�W5����
�wO�o�c˓[B��Լx�J3�V&C G�߹�K�oeZ1� D��R\�ZN��`o/� ù��C��K�_d�2g�\^$����pg���2x�"�Z��`�4q����!�_�SY�L����r�K��~�?��e3���d�B��Z��~���0�QhCv+]A��jUA��פ<�ŧ9�F���}q;j��&�E��´��e�cJ���Gῌr�*��[F�����s���&d���O�Z+F7�^s92G�E�ԫ���tcG��e�3=�1�"�� �]|%�z����8MN����G��"���	@=9|->�?���qe�b��>�5�|>Z�/�l����BoL����[*�7|�.S�df��8Բؼ�å]��e�>�8��4���� ̈� S��n�s��X٨����F��#�T\b�����HƓS�]���2�m��;���^z�	)!��_��=}K.%��Pm�+SXV���sE*T�.��_"����	�{�����=.o_#k�
����Y�.](�:E�g�5b����nr9�D��s��*��V�lNJ��M[w��O��S�<�՘c��Q��A��рD��#���+�k��\��� ��əO��P�.)�$�8��؆���e��!ԝ�q>�����O����<dQ�eSC���r�3A�����#4����nφ�!�۟j���K�6@�'�����ʇ֯6E�����K�P������+=(F�/����f�,J��RD�#���f	��M���g�
�i���zޫ��;�>ӟ���Y�]���}5,�G�)�zB5i��9,Z���!�ȣ]�]"�y���ZA��
�]��s� ՒQC@G_��)��V�S�#^M�bw~ ^l���W�y��I�8�C���!�F��*y�cD�6+t�N��n$X]i�=\,�m_3�Ep'�ԡ��L�۽K���9x6����	�������VL�D�U��⊕�/٦�N�2�y���Kꋱ⪊~5 �;��^1��Ihp�&}��PE�� ��x۸�ߣ��?�#����X;ׇ��Å}M�.]BTż�Q�<@T#�i3���\Eӭ����΃����S�㛪���Q�7-Wk��TN�O��	f#���ۧ@U\V�}���(���z���^JGc1�?�*����C�\ϣ���J��rG����i����m'صz6_ ��K����3�l&��pR�H$��S�����I�U��X�~��/�H�k�5������:k޵4KW�\[�o.���Et�?�>��=�&0c���V�ޫ�Gm�j��#wx�\�&"K������D�)P�W>��m��O����G6�~�C��h۹�� ��"�EY"��x@�*r�$ݵ��H�BtB��-s�:�-�S*pҩ�뇸&�@x�M�/�bB��L�1�"ڲ�1�cd�|���q0�L�f�l��8l:���E"h2�� F�� ���X(b���c�TJ�������/���Lo1�N�ړ2��������?��rXT��D������!"��E:Ӝ7�����T2�0@�)!ZZ����U=�j<�6v�.�)FBF�i�%���٫�zK{���b��X��P#4���6a����}M���pg)=՛ϱ��f�[��A�:�3���ɏ���~�ښ<K�M��|`8U�٥Mr����-2�iˑc�[=U
��OR1�\�ٻ�� y�L%63�ri�<�򴪏�����b�y�4�l�UP�(J��M:��mpk�TEDޛ�)�\��>��4a&ix![��}OS�}K?Ì�^���+�у�����N�dm0J��nx��Q�Q;�6%����X�O�MB�R�V����G��U��Kp�xaN��hR��,6�l�`-G�
X
�&��og� n<�� ����(b0�ޓ�*fӍݭ�`�X�@��r�٫c��<nk<��G8�l�e�+��ګ��X��L��m��a���#�o��ܿTj���1�7�,#p�:	��Q�?�'!֪}X+�\M<�v�w��cΑ�d���8����z�v�"�,��o�5/���)8�<��P4!�5e�L?�ߪ��F��߽��X9�/���)i+۝�=��L���d�#PX|	�~{c�:S�%)%��X�CU��n �2��j�� �M˛Ogrym�ߥ�}vxx�J��1�}.Ἇ%X�o.T�~�?%��<i�2��G�`�ͺ����gp���=��'���` �W^��!����`ޞ��1�[w�kģI���H��j��� �8���ĹTL����x�.z���S���N:�0 ;/�Mi0b	�������Qy��i��5 2�0�X� ��`����-q�Zz@�s!:��!��X��C͌俨��4i�vh|���%���R �LuUsU�}F��=�8�Y�Y=W�>�n� `���</LQX/�.^\�ƫlm���I�8�G����J�^Z���Ʃ��4y��0q�W�������?�L���Kr�h��U6���8UoȊ�	�ȷx ��2kM˙o�:���o)����
k��٢u����~��Z���X��g9�j�߂�󤺔o�Uu+��������/�|���X|�݌L��c��b�H˷�5�-�"��<��}eļ[�B�GH� ��E��!�t�>�0�{��Zب*h�.ҭ7�_��1<�qr2�>C�F�١ �_��d���?sue��h��*��`�6�����#~H��yI��+ߩ��c&���
f5�[>��zմ��5�}}��������賿��Q:#I��Du�9U��*BV<��Ws����c-QѹGjG�Q���"�s�t�3u�l����� ؑY\�Zk�a���O�B	�u�||�/�Dc^H��m�)�� �'yO�1R X^�N꺇�=�'a�Q�eI� 0����yr��+I'ʥ�e/�]�Ԭ&ڤ��?����s��2ɷ���ߵ���ZY|o2��X*��=�����E�Pj�՞".�Qݻ�6�X���&8�iT6�;��IT�:}���$�y��5K
B���a����������I��	����jPh�V�܆��	-����O�LV�8Շ�6�*>����#6jB\DC�� ����rO@���
�d�dq�|}*���,��)&FB���	xIw@-s"�/�d�m����<���֙��d��A��IĜ��6E'���۾��7u7q��p�Ҩ)�3ߜ<�:���G��0HH��NR)��4�=�6&nvd����u��[���(uފt��	�b���kv0Z���(�H3�,V����7x��\C}4����2�ߑv2L^bi6l���S�1����̗�hk�l�U��.r����0�����;��%�=H(�kQm�i�h��O[���U�)0k�b�AX�u��}ߌ76ݺ?z�z�mq'�FO��3�{�wi�iK>c����[v|ع��-��_�Px�YLa�ˊ
2 l�Y
]��8~�
;CB�e�%]Si�����_SP���_�r�+O%���r[	��o�#'&_V���=�\���%�S��Y1��y��S��P>o�x~Ht)1d�X���B��kG����-�̾�g���r���ڋW��8�
]U.߲�Ns?��!���e�-��}b���	"@O�M�۸=�O���N6i�M��L� �p�|��X��u��e��N�5:{B����[�\��s�PQ��w���?��pzU�G�p�xO>�m���̂w��V��雇;Ѩ�G�G�n�OY�\�� Γ���Avo {���E|ؿЇ�W�E�`�A���ޠ�%���Gz��v[�%��{S���6���	Ѭ�[��@�f b���mc9��t�p|����S�(�6]��ss��ڈp�d�8;	��V$��.ao�|��h����n���)�:X7���Krf��v��ep�}�W���6���i��-w�Z꣘�*���e��m�
o����|�ۼ�����5��c#bv�L�q�T��y�kU�V��|�-���?G������T��g�h��Ep�Z1��}���.��[����ug��[�_�=6�SL�������sBXj��K��,w�M%��y��{4�w�)T(c!rb��(d4/�������
��*l�fA���7���(�4]��j�`+җ��B�=�z]�&DkbY���1���}�>��'���F����^2��*0����|�5��J}�ş�Se3M��t0�3�w"�>�3�F#����Ȟ�,�8krRl�b
u椌�-(����i��m[>�o�g��O���� ��N<�od}!;e���~�+�r�{Iw��]�.�.R�Z�]M�C��qWj��w���E�����5�@���W���
�@Vk�u-���ܒn����д�0��"?63S{#u��T�����*��!�x�	�:}��)pt/�f�/%�4����&��A�#���<Keyd�P���E-�"�N��!�@!d���͵^t� a ,xNq���r���pѮU�ul�\}�é�^��'8��!������hf�z��Ѝ��C)C�V;H�?��'ܬU��z��C��$�o	NG>�/-�%U=�V����J��_�9��;�b�:@HX����
F/�!q 0� ��LA�7� ]ހ�wމ.!X�J��[��!Y|�b������V�[�L"�
'�C��htX43
��&������-ŦuA�����c�FT�!-��8%,���g��d�hy/�9B�R��zrO�h�5
qe�%���?�^� �[$v�`�,��8/��0W��C�����0V�'_w�8$�|q5�u!�l����H��>�޷Qӟ�����p1�or��V0��"R����%ס8k^�^E��TW�i���w�0�i��r�j=P������=�✋��q44�B��C�yQ��F��5��d�`�k-@@)۰��J���ذ��h?l$��Vu��2� �y���(�ύ�_m�%�.�G���4]Z�O{*劁�A�Z(S�oD�	͞m")��~1��ޙ�!�.�Ij!P�]/��*A@�����~A��Sj��H2��� �A�~P����apLzQ�"���)zKm>�c�P��0!�Hp+9HL�]5��K���L/�x��4x�ݎ�G�H��M�����cx��J��L���
B����LE�y���|���Y��TЈ��:oawW�½%ݑ�{7w�6w;+�E0�K��b��B�u�:!�@A�,����>ɺ@�#s'�1Sb�f�Q�*��h��>悎P��L �;��7D�F^Y����'isA��`<ţ ��"��O���a�9������B�
���N
eVez:5�C�n����K��)H62;6���5D}��6}��<a�&S�݋�e����'e*�L:�T�s0��Ō�=(�B�X(�\K�.� cWe�m���k@�-��c�� s���&����92�2���P�'=�n�3��+H���
���e����]6XC��j�h�()k��<�/.G�뷺���!��Qu`�U �4�9B>,�Yڭ�r���8�>3��	L�X�KaV]bW��_=������nf��iWKI�2�ȯk�	H����E���O�o��v�
�I�(��Muo�ZkK���O��byaG�~)lCy���縆�J�|�3(�GJ������O<�6<(ͫ3|�5�/�P��*]�Ji/=��ph��0.���t��,IM�HM��v{�R�7��}>UQ,�30n�OW	r�ږ;Ѽ�,#�CY!�����P"B3����<A-e� �"�nfZl������т^l��B�(̝k�sH��^���e�]��VH�MMmu����ʃ��1G���#��n����)�)>C��)y�C4V_�qio�v�A�^Y��Ɓ׾��y��(�9㋲��%��i����&�M�6ȭ��R�L+����ԍ0����w����`a^��a���k�G��I�����"���U^���/�Ԋ�2�G��v!Ȃ-�#?߮�[�А@�e�^�oU8Dr��Uy��_ʼ���j�Obⱨ��@�쌁�pS�M��#�V��Q��n�X^��p�iX3�h-����6�.��քT�5�Vl
S_7t�(^�����sC��a�CBx�YP�|Y�3W� ʯf԰�<�}���%(Tt�vH̫�0he��-U����5S�&��;W��L�>�E�F=J%D�,��"�(�#G�P������m��˛��|ʒfꕩ��c���G��>;|u�qV^
��I]3Q�.���?Xa���7�`9�O�8���@-&}��ݍ#�;{�(r�O�D|ߌ4�N���|���J{C^��_��_~���Q%�W+��?���
^[6�"��"��n�*%��ʾu�d��.SC(HJT�C��u�ZJ�:p����s	�l�r�mRV��SG=��k|T(w��hkfT��\*�;�m�I<���[��U���Z<nI%\?-�G��Jb�wǼ.L3�+���e�864(�~	��Xo��x��]lʃ�6J�Z��S~���j�Ly�i�oK^!yv���w�I
%t\��[�S�N&�,��N�hA
(M>RT�+�>2�x�A8�J'�G7 W��HIa.�g'��b��*�%CCj�	��8��l�+��	�=`�߷��4^��D9Ћ'�c�ղ*z?P.��w�j;�i�s��Ni,�.L�A���i2s�d�Qz�Z�34�-�0�������77K�A�k��N���D�� ���DɣA�@��ι�ag�t��@I�ّ�,�~p`q��<ȩ�
Z
��̏�UO� ��Fߡ��w�!��j?fn��18�^ ���Q0�j�Tq����4����P1I�\B&w"��eSE��k��C��o稆X}@-���}�	G�./�Y�������6����i�*�������xb%�������A�F�Df]9�G��1��c���d���'7xߦ<��:Wf� &�%�p)*�&R��k�]����$I�Z�W�-T|2�0P~��\dp �5"�ֶU��7��^5IR%�m���b��%�6�$����S�P
�Z�3W`�����u�hF^7�u� ��L�s�,������l8K׹��9�9�FrQÃΥZ ��9�rU�mo�Wv���H�Er�Q�%�۝�I�>j?O�ʣ��]�΂8���'�yS���t�:�A��{}ڭu"'&5�����<�-�j�9<���q~L�b���c>��!;;��:S,ڙ�pN����%��l�x�fJ��l7����3T:3N�,���cud�����
;
%i���qlu��ա�*��P�V ��1�=��=C�/�
zv7���ݯ���N�,�Sz�����D���s�b|���-�섶�e�i�bD��Ys�dR~5YTǙ�ΔM��&7o��h0�xH����F��}!���n��QO��ʣz�
�>�8ڍ<rU�������&���`��P���|�:���SF�&f��ז���||4�i�d�].b��;��a�ǀ%��ԑ����*��D����W"Ƚ�%W�w���H���Ғ��;�ZR�ݤ���D�F�u'�ӽ����_������+U�\��Y��&�¬6��NFl�('l��w�
�R�����hӚ�,[���-�l�@��<́齝�7���ϥ0v��SS�\��8�h\˿���;���������l��w��9��=�QUf�H׽�3#��&8�w�޻�r,�$E�Y=�2��<�j�ڔ@y�j��ui�C�|�t�0�M��aS,��A�.�tح���沸��r�˟H�a��$s���:M��ʭ)�jf��W|��~�*�<��+,��vm&�=�C\[U�Pz���*H�Kդ��ߍ1�5ì7ը��J����o�Ը��R�][�z�\/�̺��a�9-�5�}���t3��R���ٹ�G�w�_Mw[��S�N��v�R��4���V*��UCQ��@+��g�%ڈ�+�rhz��(����Ɉ�7N� �sEp�)6�cX��~�Y*t����qՒ8!q6�=�!�.�_{W��g<t6�_�K+Q����0k��{�0x(��-��ꌶY���s�z��zJH�\�%&���MO�O��M���\W��X���-�3X��umn��n|�r�N:�:!:z�D��s.���/��
��b�R`���M��$mBp�G��r��އ��%l۪�$�]{��9Pxd�t�6�Z��g��j��PMk������>C�$�-����aC(w`�Fc�I��*A�A�b���ܐ�v�_6�iT��T\ud(N�������d30	�}�(��$��n�ɧp� �ط}��4	�d��Di�T&"*܃x��h0bLK>�U�3��rA*ُ����m]u��*���$<�P��?2�M����U%`�b?J��apre�y6�p<0j-��o�T:��u���Is�s�M�5���ƻ������#m�s��}��_26ӳ�*�k^��i�׃����|�c�e��(�/wW �DW�PK����0��:=i<� *գ5�'�8��¤�U���f�%fN;!Mj���7���LK7gĻm� 
�9ug.L��� ��7u�?��5�c�UT�낼�|54�C��;e"B���6�6T����Ɵ#�,hz5��Hg��0��nmg��gp�F�]+������$�x���k�Cm��Y�s��3�2퓐d�Ǚ���|�`�k�� �p����m�"} �>���t� 2K���w���Iw�U5��do�Ӹ��-
� ��g_}?�r��"]	�n�f�g|�M1^�G:Й�4��9�,{@-���ð
5�j������HVĎr�<�밄!̈j%tK:��a�FPlf�
#Qn�e�=r��z���~�<���w܇�5p�!�E.��hXc��$���R�IR��\��
#s�ɕ�l(O>X�s�ْ�1��F6�H5Ţv`�<�`�f��@�S�ʠ(Zs{��|�H��]��10�8�s[���r�PQ́�����#�Z�����*W\�ڦ&.�к)�O����io\�hCVcM� �R�?�����ˏ�̇+̅� 8+�NV(�{;��k��J��˕�rH��3S��b�����؆��t�U�i��J�&�Q���7ñ¯� ��`��8y�j]
SL�W�_Z+me����Cw���k>N|��ۼ��
v�ԎSЖ3/V��
#������礬[rT��	OG6�)���������G��͑�"gq���}����%t�
�!eC�'�iᶎ��f��wM�l��WV��-_=�q�4��u�^\s�����wE;�b�P���$�<��׷r1������즐%C�2�!�)��=v���n�R�$��<JMB׊Z�Lz�p���mϙ&��f�k�C������H��ԛ�3��ڲ�j�g�4gJ�)a�0�A�
��J��Ε���ͷ�Y9m��"9�<�>�����"�&�0EpP�C����q����z�����{}�b���nu��3e���.����κ2��H�|�^k�i��@��Yx��f ��"(�yѹnC'��J���φs�\r.���f�V!����'F�rZ�%2׾�%����~�_�e�?���3��v>�f�m{)��v'6Gz�J���oH���\�y2X��aq0�݊�I�W2j�u�����%{���Ox���|��6v��l�_$��C�n*�c�W]���:�d��`X �����x����X޶���������z�|j�z̉ܨ0p���v �z� %�1�_,�Iw�2�2�Ql-�\�f�O!q��Bw0��D�����q����id�\6�_���;���t3�)�\@n)�����r�t�	�	�]k�euA�pQµ��N;Ef��Y�O��k�V�:4;��J�v2���f�y]���A2_�^\��ڪ{M<��L�RLT�`����qvx�o�
> 2[�٪-PRPH�=^ņ�;@�a���Z�����[ce���ȁ^��\�
*
�$�h���>+c4F	N���]1�%��������;��yC�_/3,;������!*Y������n>{!�ĠGb�s�P:�ނ-�?��6��}��3ݚвuy%vK�d$�O�JWYӜ��k<gs�f��Q��ܥ��3�0ß{�<��P2��z�����T_��8d#'����ϥ�_�)z��h�Sgv(��F�����N�fN�����To�V�uЕ� g�4˿2�=�=�;���N>�k�$+5)�)KX�v̓%e���_�Dw.�_U�G%l�;Z�i#ە�o-KC[=��T5'��%�3"�)�i^Pc����0�"���r]����B�;��3��,Q	䓦pӕ��������3��`�O����Y �>355�F�$��g�8�pO2�'^^�_a7��o��ږAA�gF��~��������޻0؋����R(k*�u�Z�hP1 �;Oc	�w�D���vU�%�i}�_��_j|���sx����E`�l�z[
^%��;\4K 6������ߠ�xK91:��Vo*�}� U'�P5�.�J� -9f�q����M���B;�|%S��j�����jDU����v}�𨧊^�wݜ�=�	�ܢQ����m��XD��#�
4�$'� Ö녋;i�����kc,��v
,����\h��|�_k�r�y�zbd��X'�P��_��O]����f��(}���s���y�@Tg��mUt1r���Re6�F��vZo���	�G6���ŧ��KGu	�ؐ
'ó%�Ş��� �7����.8D�Е�9�A�X��k��ʹߝ�4z!��k�j��������1Jͦ�YoĞa�	j�@���L�
%_�yH�Op�ԣ��V.�p8�JRo!$/�uƽ�=��<�d��c��U6�#�c�DY�@���L%"^fk��y��T+M��^�cE��@;��Ք{���$��ַ8�J��ě��Sh��/�)��U]w2�ܙ�/[ud�y�Q�Y�T��H�}&	��FԆjDaySs�J�|ůe���� ��S���K��x>qm��pw�����W��Eգ�M��Ŝ���J/2��d�t�IӾM�hd���/��@�zk�_�5�v�E(���Ȕn��ٮJ���p�9�"�����T��I��P|�(9�Cd��
��M�b��ʂ�Ĝjɥ)j`H��v��,�]?f1q[��w*��A�E�ny
Xn4�L�Gp�;5�3
-o��ƞ���!?-c#��'��'x�oIb ��q�_�y2��:���5O�1�mz�;ҕ׌��$r���x���n℅���<�+�ֺ5�Xd�4N�s���� \��*P��O�
�[oa|99"\�`9M����q˴)6�)�U�E}�b�ӜK��� [��i�+c3m\T�kB^�d�I�ϳ�>\�T�`�~MR�\>V
��\(��^7�+�h�_L��%Ρ�:�;�����"@1�׈�@9�T��.�����.y�ϰ���E^�Fh$ݓ�{����ǇF'�d`�ײ����m�L�kl����ê�C����b�t��ӷ{�ܗ��zV��+̜�Ç-Gѕ�{���:+ː#&H�]�j|aR�mQ`������0�ʥ��$�I�o���TY�bL��T݈��2��hR�L6ʇ��+�gn�ٌ�0Pb������އ8�v�M���i�}`hrm���ʯ������fMi���� ����P�p��s�j�:6�2���.�4���u�P?�?±2 @u����頇�^Q׌��F�E&e4����a�����dD��*Jy����Z�X�j� ������bٵd�Y��H�� (��H���D���3ĶV?ʶ��l����E�p��G7��({��H�����n<Lڎ��Dٿ�0L�A�W�2X��HGN�����\��(��>Z,���ۀ<`i`F��S�+x�n��<����a��y!(��U�.��Ak�ƫb�a��\ݰa�>i#M��z˽���N���M�f�rDo,��/V���%ƞ��?�s�2���!vOs+uLI9���@j��*^3J��v����}��-�>��_���U�H�-!�#�o�]B�ߛ�WG߷F~ ���u�&g|�K����U���qČ�D:�#���a�8,C�A7��g{����b���%ԟ/%{.���N�H]mR����x�,1�)��f��y�3�}s�B��?�,L�P���Ҝ Zg�� `�`�m���ݫ
7� X�5��<R�w���?`(�seiD@w9�,4Ã5j���U��O�Ja�y���H
w��7,߼�i(��S�3��0�f��u���x��ei�&��OH�RӔZ�4ǃ���L��ML�<������v�ʹ&��ݝ׋�w����j�a����7{cƝ�[<�Zׄ'�q\�2���5Z��1�� ȜS<A ����?��wy,,��r��(���)�1��y@f���[�!�4��ǝ�TY	�:�Yt���&n�J`x�rkኇA|��/^M����^��ID`�x8��cmB�LeKp^�0�M���G�$yF6W�sz�V_��� �`N���=(�'Z�]O$<��%E-�ȟ���O��7=q'�/5V���ّ����i�Y�ُF)ٟe�S"j×2��h�aw���1u$V����	�&�rT�U�L[��3q)�:d�bi��^~𭬢ӖI���V��u�'������-f3�)+�k��m�&�>�H��cނ4�Uz ә��w[f���-���˽e��Q)�t\�)�k��M0G�g�x�|o�d���!����W�t�b���1�p�~*��{�w8K���蝄AHq�G��g��R5���}?�XE��L��|�X�߁Ī�,����I�%�N��g�n�d�M��7B�b��~�7+�{��ؗk��\�W[n��1�����V�ê�PK;/%M���q������Z�]cwlb[<�F&�f��=�B�V��J�� �_�^��9H��ay��B�� /�O�֩4�ת_h;Y�,N�闁1�/��| q��.���?GL����2y���^Cs���5ѷ`Z��[��4��bDl׸�x�
F5j�'-� ��~�&����=?��K��I���vMLr|��h4�n-Ǆ `n�䗼?�q��}
�01X���jMV�,-0}�6��s9G0b�g�)Ds��bI�F���g�S�vq���8dR�g!�f�N2��`��:U���:����k�4IN�����؇��� z�'���w���&TF�>_38�ܺym��0����ּ����$�[����$��|w�jY�3�ɍ����i�5(zĽD	X@��$4�_D��=_��۶����PÅ�"���oF�Yˠ��U��`H*��҄�n/�3L�P� ��K	P<Vyӝ�&�`�����ޮi��a��ᇋ����`G"��}����X��#J ���$�tG� 7{"�`8�]���-� �*�č��ϮFƷ_�{��J?½�9;�&q�G�
�?]�!�?Z>�k>W�a�4���oe���fB��oV�3wC�%'�%�Z�x�D�d�-:efߵ^��\�͡�uP�qjͥ����ThS?Z�d���o�����ˁ�S��P�,ӡ���&�h|��}������lx�%޶:S�/�R<�~��_�������8��Ϊ%M8e]�w�=d ��5��. x��dX�u�qV���%s^m�L������	���<�+^etB���Z���1��:���Ů;,�8�ZH���QH��c������2ĆU~�4����H�,���"��6���%}�)�U���<pO_m"|�~ߛ����g��ă�Ѫ(~P����s@ʋ%N�C%UR���%�J�:L�U���U�j��&���Oy�A)`��0��{xP�|�R�R���+�.z�X&�W��c.�f�wL�����!��-�����_+oFv��$�<�#[dD��@ʒ������p�79��t�p�S��ڵeC����y:���������N�~j���jo��ƺ���k�NI� ��6�����(��^�n�)OvJ�OG���nRBR?ӟ?9S��y��k�������E]�"`v-�~}
mE�A�y-D�Sv�"TFs�� ����0���c�C���ANQ��������r�>ÖD�pÛ�>��+��f�A[��ӬC~�O%-=a��V�50�k{&�LЬ�RM�������h�P�P�l��qd���Ln{%eB��_���m<�U@�Z�0Y��ﱓ��(��\�D�����,��I�L+	R]��K��3��&֯�����%yY�Q���<�|A?Ď&,8M��7K�^f/.~R�z;�$�UX��z�{w��04]1,�c�8��Jf�B��jr�b�*���~���jl2J������Y7G�Lx���Y洓^`�������b�yp�A�̪>ŕ�A*�i1Y�������*c������^Uo��l���CS͛���Qb�4m3���3�=l��p�W�s�����Z���drU���be��R7g�[��x;Z�e&�+�G4�-@�vf�y��������#�!���k��ki&�<�yW%k��K�4Pn�(s��Y4B�6��$w�x����Y�측R�����	&�t
�S�[�����
O_��'0 �ck���);����ƺ�b�M{���s�uT��fja�s_t�j����v_j�!1��`�&�lyC�Mu�J���'���%�0�Z�e��}i�;�	�7�n��CT��f
W8�OZ0�M�}Y�luXK���K�t��I�Q%�W��y.��h�I�^�T�B|�ǭ�*|R�sT�W{� �ZO�2փ�ڹI�v-�����M�c���붋��(��p ��)��������+,���V�,ٜlAQ�=4=�Z��ߵ��iD_N��i�YP�aΏ�B���g�GiP����_���A�M�ّ��t��1p59�_+	�EN�ߴg-� 6-��k�o�#�U�� ��#�+{�K��ۅ+�d�]�]°U�Y"�d)*b���f",g�t��ɛ1�8��ۯ��3tT�K�n8g�6�I�i��C�TkEhj^H7�ڇo�Jr�y�r�-2]��1��$u������l��8HƔ >�}�~�Y�C�/v��P>�W�0#�?����O�!��!}���8�!�Lo�C�#C��vl02�rj�b�R��A��q}��`���%l���ق"�G�*����a�CZI�W0���[fGqw2���Ve��$�"��� 2�n�Y�qz�^ҽ�h᪪�O��nt��1^��Ą�e�<�`�L��͡����|��6�1���M��H����\X�6�o��y!o�i~����Â�>�ߙ�%�Ds��9!�7�!H�q���x�o�<2���%���H=t����C�Qu�ݥ��	l�*$q1p�������oA[W"u>eTCR�k@[�^�43gn�fl�zvN`�#*��P|
X�y��l�DҜ��7<��x72�5H��>����X]�����ћ�n��>n�]��K� |��e-��l�?nM������>��3����/� �~E�5�e4���K������ZDF:��&�E���4�F0pj�ל��C:[�H�İ����پ�݉��J3$E�iD�nސ�����%�ܷ-��:U/� EA��[�E_#\{�Yo����g�e�I-���w#�^�̉��CJ�{1�Y?$���⢥]��/(� m_�3�`g������$H��~�d���_w�ҷ��]��5U�ұ��W��a׽N�ً��6b3�/q�Nm2�0�&�6�ͮ٬���"�w�30�0��괏�
�d��!&,܋�X�s^�΂�&���7Á�S�fv�&���H���K�0?��E��uG@H���r�@@U�T�%��v�-�Vj�ƶSh�ͱQ��A�Q��g��V��S��3�\Ojc\�*��1mOQ��.qF }�0k���ڿ�N���:= W�aG��&�ph���R�@���Nag��0�ӂ����2J��J~/cH]��d��UCd�vĴ6�g�\������������,�I������3�
{xܦ�hۘ���C�*��5V�P0�8H�\�))��2�]�?Da�k�w��
u#��I�FA��ln2�~��gV�`őWB͝�tf�0���tU<B�	=�m�D���`�pzM=W���,ky�˜w�|�N��x#�gb��B�-k��}�C6�@�6;LǂB���RI���t���e�х��Ou�'ٰHu�4�2Ad< ��X`�r��e�!������Š��<��	�\w*�z��P�Д�գ���b9�,Ǐ5�J 3[�����!��(+凋�	sh��Gs��z��ܛW�|Ō�����B��]��F�p�6��� �.hvj�n�v�H��R�~��
����k���+�ҿ�%�j!v�����Hty~AC�K���ardy�3� �Q�^}���$=����P�	C����Q�G��I�9��]�@�}�R�;CX*��Qzm����=��ـ��Wͧ�^oׂ#Wۯ�iS_=|�w����.�:�c�w��~���V}�{ɲ�+j��#�6<�mp��М5׬�#���j�CA�R�͏��v樗*�|���|�WB>rTM��$G�Ij��������:8HÎ7��gʵT&����($�^�2����2�"��>�c�p�9qQ�Qia6���=�U%49�������)�HU®dG%��J�S °-�#�ӗo�O�$7լ��j;Mq>7N�ĝ�:o�k^�"j�{��_�����q%�_<�0G9*�6�xQ�i6&Ai>����N����� ���6�F� ƾ<9�c�i
��p�~׭+�nC"h#_�RsčZ=�*�h���A��TO!��넁	�V���7��_w�#��fOV��W1Ȧ�]���vB&Q�\,�kܮ�Pa�ݿ�������N�T�8��#�f��C��?9���,��׈����v*A������^�qj� /�ƾ-�\H�sN0�C3�����Pbr������ђUG ����L������]G2�x|,���9@4u�G���2�O�����|����t�����&iXE��%�K=���SYq��w Q�7K��]��#�e#��0�S5"ÕbK��P�A1��ϷKR��PX��ʇҺ��C'qlT��_��\rE�Bx���}U���/Q�%o5"Td±=~���w�+g �'Hz��Kmn8!���l�q4f'$��",H��Ei��6������U\�E˛�N���ÚˊK�h�_���C�]P�M����C�(���Z?e̅�7��d���+��Q�13��w�*���&���c��u�ʚ'��帶jK�Ε�e;���@O���U�
���|�l��;�Y�R�tX�:���hv Z"��ѧ "P�z��90���<����ᥟ�9��d��3E�1=yQ(r����R�Ui/��n��Α�c��)�S���~:G�^��{Մ�e��md�ՙ?(�o�,�!_dN4 �4���E�߫�/v�y|	BŦ�d�d�S�+e� 'S�5<^�q�������=-�Ny�&��J4j\kr@k�Y��\���j�Xa�
H��~�%@c	�2�`���J\-`&���F)_"-9sC����Y�xH}w��[��+��;����֭�:ڷG�9cZwy�C��^�U6��؊n��ʥ�G��@�c��!�N7�A��]x.����T�c��i�k�y���E/��4A8]͉B��W*Q�`��v$;��a�2���R��/{��9z�y�L��\�h�B�h��W��_��2��6�m�O�:ʫ���$>������Z���W���ʼ�����/���`��Z�B��	����˜��wbeBB��h��F�)E�i��~c�7���yz�0� cÅx�C�G�/70l��g����[��z�0JdL ��[q�z��lg��������wZ��y7R\%ҩ'W�ޛq�v�C�,x�%�Es�������&3@>	l�aמ�'�X�jL�
l��-��N�N������U�+� ��ԇ 4#����# �Ќk�XC�X{k�Q�hk�6[]�ZӱS���_!�&��f	GK�9����,9,���i.PK���+c��+���$0^�i�_��>b��{�(L�0�ۯH����c�X�����a(S%�� =��,+��5�� R�#U����?,G���!�GK m��z�(�q���!�PQ�֤D:���v*Y�}�ӽi?�	A��# ���������*��_������V��1�3z��ݒ��-l��=w+"��\ ��T��#w�2˔w��'ue֑�UOq��k�:�]J��%��8��o)J��1>�����p�@I"z$/r��jED��o���3� V�U��=�'�v*��H+�߉4	��ba���)fɄ#kR�����	�H9h�~��S�U�����lH��Wۢv]��8�"����1NJ#;(Ѧ�})�<������sqB6JJN_�HW�I�O)�Ħ�;�[NL۳��b��G�t��m���}�W�	c·BF)�&�a%�M�b�ڻ ys�O�X�9��� �kT��*V��'f�;:��ID{6� �mhfނh	8G��R�q���V��`���P��0�`�Z�WOHҖy`[��������P�+Dr'�}�Wv4��e����H«�Ի��=�J�v�������Fl�������im�F(H��3���D�~���/9��_��z�ָ�����53�N
�$����}��@<,��Ud-s.�����T�*s���^Á�����,J-W�{��p�#z�(�5hYU�^�k��pL=�'}�[�����{��bN*���&*�y�*s�Q�x�r�ĸ�H�X��2(%%W#��H�K��FT�.�g��A<8Ļ����$�գ��mPa��a�5���Q�d���ɘ%��3��ȯ��f7����:ي��)A��@����;�\��*�0p��N�bUV>X��M�M�{�pOF��5'�O:��'�ߪ�p���r#�녬��A̻�n_�8��Z��4�q�?u 1�#v��_�ء(Pʩ��v����^�%��#ݜ.�h&$f_b� @*�m�e�`f���$ڠ��(pc!��k�o�m��!��G1xUL]f�i=�K��(��� �0mx(����g���'�p����bV����c	@���3�:�p�n+˜�teޥ"�6�ٍ��9� �m/��~�s@�:g� D:>��o�:"|�I�gA�ާ�����a�F;Nr��{v�γ�)6�q��	"��M�YyI_w^5aR��rO-E��@S�6z�J#��5�����XIG��*��v�\�Mk1l]�p���n���Y�5��l�|5t���C��z����Ht���]�0�^ү��$�"0�� [���z����1
$+����/C#�4�6�q
͵���|1892������p�����v}K��:p�Dc��Y[U��6rI��8=񢞳�W0W}��؃�0�{y+ۗ�#Dj��"� �#1+�@Dvl��.�e�u�:	�GW��m���m���BA��3_������};^0�,>$����mC��}OA/ݬvG�9o|^w�FR*�2��=T�2�5��E����mu���OO)��֜��ĩ���ҿ���a$(���P����Իţ��
y��0�嗜{�q�:��dZ1p5����-��!��?���i��e�{��"��v^f@�*��M>ǵ�n*�y����&dv�o�� @'YWs8�=�,FTu�%�Nw�u;�o�i'W:K�` ���ԯ͢��W8"�!_����W@��� [�l=A�Į��]�h{�Q��C@�����5E�� g+p�~9Y�z1h�5��*��O��j�$@K��'%�0�=۫�r/�: �_? lۋ����[��n\��]o�^Xo���t���'�NS﨓��Zڗ
zY���zM;z��X��}�Y�oc�(��9�,ɍ�u\����C�o����Bf�#�8�ǂ�k�,��jw� �p�Abw��8(H�E>�r�د��_6�f�:a��ۧ���9�xg0U�U����B~�c�f�c)$IF��/���Fmm��D��z�-��ê�f�J��W�1S�֟Ҹ+��]��5d&�O���|2/"�=r��z�Me�|�W3���������y���Z64қ�`1LR��Z(�����/��ÕZ�D����lb�R/��bX0�mr��TG�I����98���c����e����7�Y/i,NcJw�L������C�"���ҳz�t�)�ط7*��PC��}l9�L=��D���V��I�g�^��*�Q��Cw(�"�4���"��>�c �iw������1�:�un���� .ʸR�����5�CKܬ�@���k��_����i�8��q��>�8����F�W��>�:se�q��Z��:�XW�?ӣw ��B3�6���$X<�?�3���X��M���U;Ѕ�$U\j�ʹ%�'��Rr28�敋0�u��'a��c�@�)�a=�=56+�@g>lV�U��h�r� ����Xwm�����&�rj�$x����獡���=D�	l�u�D�F����6PQ���"��AQ5���0 ���TBb�_ŪGޢ)2�X���g'!}.��<��BU-���Kf���t�	m�kg{�Ǣd�W�:��Kx|_�Wz�?~��O�|�Ed	�y䫖u3RY+O;��{F�o�!�ڌ�K�'�d����c���*_�8��C�� �ʦ��r�O��G6��>���ڌU��-Y9��QΖ�^�*��T爺���Kcڀ���ߩ��S d_��'M
��{������!#���B���ڟ&d@�{-")�X5K�������}�z@�0ء`�c{�����sW���y�V�&KNt&YC
�J�'ӀLW����	4����Z	���x԰��~�F�)���zq�;��')�fw��x܀R��*8��3�U��1L`kOĞ���z���iD�f�د�F��\?��¬%�@wr"Q-A
��	�)Ӫ�6���M�3�0E&���ݪav���	�Du�K^��.\ P!A�Υ��]񓥔����Cs^��&�Ʈl�P,N�|�({ 0�{�5�k�}�:��g����.�-�V���Ę�᧨|q����_��
�l�j|��3��\=p��z��E݅�~��~:�TQ�(��J�K]���(d�;�\�c���(9��bX�'k5ȸ�T�T�uĽO ߃6QV�
��8��c͒ [V�9�k.�v���W�YZO �z��y�C�.9֣�P/�p�L"
��&�U���?�sm�.[��&�f�|�j� �:���c0�����0�Ȫ�s�`5Ț���m�f��Po#C�4p�@�s�=��M���t��{�^Q�r���߱�q��J��M�6i]�w�`N͢bͽ�5Ad��ג�y.�i�{Y�(��My���g�4xf�[�ç�]*8yT����g�����>��
-x=��r=�'�,l<�K�^��� �}jH�g��B��W��ww���ǐ�V�T��zY�O �u�2���z��7[�#�!� �-�?����#�k���=�)(�g�`�7��k��C*��C�+�r�gC�ħݳ��%�@��]g��go[����\�� 71����R�e�=��Z�T�̬*�Խ�͞����^�!#��0n�`]�zF�V���X����}��|����dd6���P|��fô�'-*	L�V��޶���} �Q;���:O��ŕ���#Q+8��N�m|g���F���2�lVS�N<	�h��5q�WAmv
0����<���+#%�#TGCĹ�a�c'ИA0��!��(�ʢ��/�6FjƕHL`T4����,����Qv� F��V`[�b�����}�򿘪[�}u� U窧� .��;zl�:�o���qS��� .;c:/� ��g��[�i�q����5��:��@dhA�j�Yk)o�`���i�M ���6e9v$}!*��F���}��,Q~乧���{�ubP{�yF�Ud�E�����NGa����*��=Z��.H���Т4�n�J�s�o'��|w����̝dz����a�8�oy�\��j��*bX�y]Hs��"��n}k_P��d��(`C��D(�y	��'�X�����j$3��G�@��"�*C)v��{�hПK���!0���	iSR���x~H�i��M-�y�I���M�0m�%oYl��ۢ	�*H�{�X`uX�K�*..�~�f��pO�շ�X3�~����5�Ķ�P#Ѿo<a�gsD���$�;���k��5gF"?���z��b�.�^r��(��E�'&� ����a}rC�a�9��G�*'>��>",�������b��o���sL�p;�lz���j 1��M��F�D]�������~?Y�W��vТ1�<�u7�{���V���Hȷ��<p/����0N<�JO��'*�w{R���1�+?��Z����N!m��oF�J��'l&���CVf��6ldʬ�߃T�7Y�ݬ�'��`�#o1p�69��O��*d�z�'ޚ�h$�B�~4�a��#Y�+>S���Yg�-cU�2�>��<��p>�Q}��^���O���1qrr��X�tfZ 9Q�Z]w���0�|��;��Tq�o�٤�S*B�/��6�dcn�E�]�7y�茮)//� {P���׿^�&�؅=��o��"�HyV���o��7�Gg�^&, v$��n�a����m]�6�ҭ?�j��;/8����雖Yt��c�U�\����]��O*�ۛYz��:K�ĲT\Dܰ���'Tg ��)�u;�A�R3�"
Z��Jn)h�5�F��K�9P �I�0��ܪ���}�����.5�v#h?�|�~�����w7o;:u�$)��o#a�]A[e��7�I/�O� c��ت	�YB*䚂��Z��\{����n�D�������h +��M�`;��L$ۯk�/;��y�?����$T�
�~��Ϟ ���y�x���d����^/�i e�?^#@!�h͹^�%ݫ�q�(ၐ��#wt�F��v�Ñ��}�UդK�(�,tW�<V���όC|�9Z�߹^X
Y|LA�`�r�&F�GPk���J�*���GGu���6�~�9ZVu~��W �(��|��� �Z�������D2���?gJȾ�+2{`���i��O�,��d"�u�k;�gT/6|�&�*�	�^�=����$���>Q{�(�`�Ǔ��_� ����+�^���[z���Y�	��l�q�i��V`M�DsaC���L}���LXI-����%���eD�+�,K�j��B>w�q�_jGɌ�F3�����n�̓E����㞎>6i{���L��*`���UҌ��h=L��vz����PkCn9�z�~��c%r~��Z���=�
�����E"٢��|�?)x:�Oa*σײ���~rf��%4 0���C�\aP�
�K�Q�y��!ҥ*�=.��P���UR0E2��4&i��WtΒ�����ρƑsγ�193�$5o+i�}�,�'�^�A��D��J gv�۞>���j�c��tѮ�)�"�O�X!㗬�b��d[�Z�X֋�ZT�'���70Y�$*#�@'���f(��pyE"��׻ͯ�_�D�N������b�d��NE�A�.�u�P$�N��Ї�t�ܝ�B��j��Me��g3�����B8�v*}�2�`�ǔ����R�u�*yq)��?�V�,uU]x��S��,k���*ԩ���4t�w6����FGe%\��}����ј�F��t�#��7���MLc�y�hUR�9@cv� ���Y�!����3k�e�M�=�u+e@0�F[ŜE#�.�WRuz��hB�±�b���B3T�@�\��?�<��J6;�T�������u{f�,��Pe3�;�Чi8��Mt-H"��D�m��*M�Ѩ�,A?g�!����)�eeH��xoz�͎��le���5HK幸�^�jτ���+Kp�Dbq���q�B5䩾� m 4C.�/ܓW�U�p@��S�X��������)�.��y
��/ϖ�(M ��S;� rHU���l f�_��x.�^� 0ΏҊcV1K��w��;�-9�L@�|�]�SYxL�aB��[c"'��*�x���$u���~ۀ�w:OJ\��f���Q�֩z���h�?E����1����SN�	:�`$�ۺH(�����/�?��+<��n���v!��$D�Ԭ��$�Ӫו�����L������,��=OHz~��Z��[p�Er�ǘ�y͆��]��A^l1.-���W���i4β�Hf��Q���71�7������J
V�jt��s�[�*sZ&�k-���Xl*�C��Eo�oNv��/)�Bc�V@��Y�"d� T��"���a��ܙ!^X���-m�}��-�~e[?��WE3��gId��4$���H���F��qK�~�GT�K��p�oQ������tq������Gl��Z�ć��^�mIР������6��+��ؙ�nS� 1��H�&Q��=GxU�@�{/_KC����-��s�;c� �@`|�h�+ʊ^e5!-j�L�F�P1jP��ջ������(�3�i���"��?"��)g��������D��Ǭ�^�Gh���1n A�Dy��H���}ddҪ�|?�0f�ӕ+bbmT;���h1W8A��|AɋF�{�Fo����M��/��GK�T�*к�opg�/u���0.����F7�P�Ɨ�����^Yq��T�ba�H���Y���������=�y($SS��o3�M�Zw�Οx#$)������lD�l��Oҗ�s����e��� T*e���qz_F�2���������9��'|��A��i�b��&������� �C��Pg�L���qy��_���ߙ�� �.��|}%���`̡�5y�}n���؎��Q>����˼�z痌*��ox}�(%�7S�ѽC��Ge�����Is�q���Q�h�p\:�L�#&�Pᶟ��x�Kz]���v��f�養�p�~��rQD���wrE��$;��r߹��aE��ü �i�0B�@�d��~E�b9O���t��Ӹ�G�;��ï��f��؉�f
�z�����g�p�.�i��U�*SB�f�B���FK*1�]�֒��ȴօ[Zy�D@�����$%����MY�8�^,��N�?�Wm@���]��G�[cp����R�2|���r5%�&��[Y�gS�v��i��W*�g��,�Vܠ���n
hWҧ�Mʬ��k��IU���A�A#�U5j�����~iҷ��I�����x�CÍ���
��Rӑ�Sf?�DSe��j��>��$�����-50�ԩ��Be���AL���� iy���n�h1�.q�J�W'�[� O��5*7�ф��󍼣+��6LͰ�r�"�^�a�>�e֍�E d������՟��O�Z�0��T�.\J�ά@nIѮkJ���!*�_]�ȉn!Y}v�����.�3��"�]�6糞�o�:�����W����jڍ2���m5g/��
@H*�!2{�L�� ��t]��He6��}��5��:6w�O#�R�a.-6�����AH㆑�
���`J������L��	����KP�*��;L�����$����+<�efxp.���4��	���a�_)�'qA�����)/DB�{��X����"[L�r+���kj�3�4>���8�AFt��N%\M/��C7Ͳ_	Y�������]4p�м4%��A�H@���M�r���tF�!0j�ԏ�Ï�g�`�E����W��Jf��7B�m���C���9*6b�	*��x`������ǿ�|p_�sR�Ӑ�F��$�ihˁ�����w�|Tq0�jl-6
ӫ��x,x�X��r'@1��:��Luo�A+�pxzp:N�V�q5���븿����7���:*T���K�m]�]��:���'�DITe>�'?H)������#��h$���$:y̥d�K(mi Tm;�Q��5Y{����4*J�y1"|�3�op��Bv�{Z������`(�<�6��e:߃��������/���!L���Ӆ#��w�z��D���26L��2�����d��n}�w�l�~U�j��Ne��k2���ǿ/��%J�:����KU�CS���.}<�vR�2{��Y��8y�<�O_#���(�P��x�L!�|R0��Ȋ��B�(Q�� ����QC����
7l'Y�lX�lw��V�Ϟ�:���o�e�t9��Y�jpr��f�W���o�{�H�/�����Bz4�:ϔ˥�o?��"�꿣�(M#�o�i������ThF���{S4-_��b�W�".��u���i����}��p'L���u�����=z���~fQ�;y%:9.+�q�@����GX߫���Il9&��B^s�B�P�C�AĽ}��]�K�t��+*W���xMnZ+T���"a�|�WO��z��ؙʊ73S����#�%�J9��9���\�0��{�:�¿�B���l��4m�+a�M��,ʯm��v�qs���P���g���,%5G�V҉�}����*��2<�n�Pi�o�L\<	��1�ˈ/�<˗�9HV�α�bŬ�8��%��J�KH���_��r}��ߌu�����:����|�*^���+�Q���{yIQ]FdE� uX�#-�T��r�*k���6sws)�(Z��NP��Ɏ #9M3#���}s4�xWY7Cz�q�'=e@\�'V�T��q{wp���~^h�ה�����m��������\�*ٿ�#�!��c��m�.�r�X�]M�%��地��ű7y=/�n{oD�a��ضx=u�4$J��.L�>�#�u�����i�A����s���t'�v����"����h0H���K��^3��R��+(q�/f��v�Ӻ7"��]�Ag�,ԣ��da�	�Q)��9�d��A�P�4��v6G���IǵsE�T2�@?��~�c �X�So�2�iAܓ�B�(c*��\a.�\{p�d��(��+��2����R�5r{�����q�H��wt0Ɉ��|P:L��7]�(�B(��[���d����T�Y�#`�:���hdk*�S%�v/�09F�S�D�j�#��itOr^��J��)з��x\��oZr2���j��sa�fk�`+%�G�{G\K��԰B��Ҿ���&�^\b5�3󷈉���U�"	b� L.G�?A&�/>J�FX��6�C��<U�E#�q�\�a�U�9�s�fnGy�s�o����S� r�\��o��@2�.h���P�Lx�9Z_1��Kf���=��Y ��qn,�z(�u
\� j=�����%]�Uz%mY�m�dr�7�<�Wh9N�Xu��km��C�>߶���A>�͊��(� ��9���O6�#�_�Y0��j�h�I�g.��ڍU���d��9!y co�U�hB�!mت�����R���h9�㛺�;���NM��X���h��sLoG�X�GR�B�E���2�6����+oYMy#�}A"�Fi+�ij]8-�#��ܼ��.� ��q�B��Ȋ1���,�簂糣�.�yX|�|�D��a1���� �qز��L`���.���=ځ8&JoM�i;���9����7ʌCƒ�Ȋ
Х�L����
]V$U�C�<@��F�i����#`���2�GT7uQмx���4�R�l���%���`��Z�H�>��v���׫"8�5=|k�`2��n
�߁�=E8���H5�S���I��v�ޑ��X�α�J�1p��ߌґ��06��bg�?1I�qBs��ۤ��K'��y�K��C�D�F����X����Nx��'�v�jl��5��a�!ʟ��VW���e�\�3p0#�)5peE��䲛��.��f��� =}BqrH�P�O�qm�l�>X!�I�R�
��.�"���+��>��6�$n`*����� >�4I����ԁ�i�A$N���޼��i�s�YE�Vzu��Gy�������s��2Ub�,� ��@�N+ʫ�^:���٪�C�b�;L?����৐g���`^'��测JpCB�Y�M+48q#�b]v_Q�ۿ�G>����'�  v�������P��a:F��^T�--�6��fЛ@�>5y܇-�}z����]$6����ݹ;��]�^Ph��{w�s;�V[���Q=���O&fPC�8K��5��
�
덽q"D$E{rUP�[���:RR���s�y8�[�!��I>�?.a: �P|+
��jo�J]�AsD�N���M�<�� ��'gzѠ��ͯ?�|�Q�*�0��Z�>�ST�a��.��+�0Ek�2���^�1�E>����|�w���!n�B����e�0��j9��b�T�i(����l�Po�l�����[X��23��n�	����פ ?u��0��2���=#�����&����̈́W������:4�3�#7e�1��梈�O|���J����{pA7a<IF��C��$ƋðjZ��[�MeIbG���豔1RM'NGL�D�����>���Nx;���s������������c'�_���U|�جf$�)a������߹+`�ag����N�SS~��d� e"hA�O��hd\����.�x%S�|�y��Zl_�s#ڌVbY���Y��uq���G��~s�A��
Est��Z�yvlA.���RB����>�XF.?�D�r��v��)]0Ȗ]�	�,����LH1�K�� p�h�M��t��5�1���X���ӝ�{�:�����h^6z�.��)�� �zY��A�f*�R�]�ti�f�C��L�
f����1�ޓ5!����V�!�΀������{J��y�^��J1��Td�>�� �`D&Nf�b��pT #�gҦ��_ Nzo���LU�wn ^�v0�yo�4����A_�M+^7���AN?���	<`��CD|�����'�ΚL�A�طBZ	�S&�u.=(�[1�a���]�2��Y�)�S�Y[�9�%ݖ��5���Iu�&�sB�ǉӱ�2��O)is��ˊwL���os��Ö�46k���>MS���ao�ߓ��"�G����E������,�b_/[�$Vt��~�o��s�;$A0�����3Ġu�Z�1�Ǐ+ �"���+x<M��6�Pb2�V	����:����7SD΃^��H�uqT2�iC��دG�_M�t>]�Ǻ�]�ĩ��6�7
2ݮ������> �
�I7�_�����Ό�yr�>�l�#4����ekD�)��t����;|��*����
�Q����I#�����_�/��W#4e������y���?f;Y&'��$y�c���?
�O�@��[��>�]�ɰ�
] _^�������T�Tk0(��Oh�T���F����M�AW���T���*]�R��uk9�,��8�  W<�\��Ӏ;�d% �~ErY���������Cg븉쾲y��,T�ohC���������|EZ&�~&F���n2	�1C�$ՀwYO�0y3.Y_�S��*���̭�{T�'�4"��:@ԂX�A+{0�; UPD�Q$�����(/*�R񆛜!]p�`��%}���F�cC�w�=��3�F��U�t���z�i�H����4'I���"+Wb�����s�k�h..��X�`�?�����hS@7�2Cͯ�o���%�ʐ��4�L���DB��~�c���E�-?��7?>6`,��l��|�aT�1MbT[�6,���8IM��%��e��⧘�2�7��HXl��º���U�h�t�f%��h��9r@�X��W�cEʢ�%��j�)���=�EOua�,�߸+�� ���MN[�6�/&���Op��"��E7>���!��eoa��ۘ�p���D$�P������,����6z�Yn4D�U�rj�da�X�6|2����d�"
M����00��������캃�Wm[q'֝w~,(Uy]���g$X���c����*���W\�#���\�;dMOg]b%a&�W��?�� �U�4�Oq���W����Z�z��oG*("�v�ag�P͝�_`e^X����ҁ��Y�y��~;^a�-�c�:Bn�0�+��9��X�(�9�ddI��f�S@�<�p6������-^��3\G+1t7'�(��<���!��H�<M��cv�O��V��!cD�S�)���o�)�޳��{ ���������ūu�4�����#��-.���K	u���]מ�~�2 �as�=2�*��%S�q�(�SA�Z�%}0�x�J��W�#���Ņ��1�b�����7�����Ìag%�v�ŧ6���Vkf�E�XY$�6�^�bDG/2Q��L^W��&m��3��S;��Ω: �����lYk��T͵��+`aU&��}Wb/��A�$V�z�ꅒ��� S�*��ý6�a�-ٗ[e�X�n���e�	����R)h�v��_��_d����.`|���#]"p��f�k�Ht/�Ħ�J_�Z�ʪ���c�-�y�k-�-���_����Z�-w	d��HaO�N��� 1h�W�i��R�f���~�𴰓�U�q�C{l������=�ڂL&�`(������FB��>�[eVd�nu�]Z�MN8�Eg�2�!��2,�Y�N`��gSc43�R�ˣ`;��?�� X`U��<`�T'��
�)��$���ޫ��:.�>%�oWm�"�>�(�/�{�1}4���������P)"ʾ�<��4
��p�t�� S�4�4���M�N*Yg`�R��?�3���쒚�Я��|��B�SٛMM�iyh�\�z�
�&�T�+	�Nga��pUtG]��6j�Sً�Ֆ<����P�n�(@E� I�>���J�T�6�����S3�2p�p"�XDw���9�Op�x�؍�'dۜ0�O.n���D�mJ�K̨Q�Q��&��YCq�{M�K��#�����M�,���j;�Dˠj�p��Ha�V�@yS�"$�DʏS�s�\�uJ-
��r�gD$�J�?��Z������m&���m��|�������1ɖ%Jc��kS� >*/�|3�����3=FG7tf)�&�	�PR���3���^����*&@Ev�lw��ktp�GZ�=�h�y,��f${Wv����X�Z���iM�S�st�F�S���eӓkW[�Q
�6���gOLX4��%��69O����8̇>.]%�Ƥ>�K�y*q����T-��b�?9�0M���ͷj&�6tіU	oC�
j�s��G��~F�R��!Zu�8��"��t� #(U1�Q��K_���!���ؐJ*uz���/���"K�ag,&�l�~|_q��{[�h�"D��!Q�0����(�-���Dg����˖;q�ޟ0��(��e��K%v��J}܃c�]��5����
i'��Aa��[e�S���b�J�7�Y,�����so�`��$�Ez�{��Y"X�6lټ��~���>C��X��ڨ�RC�Oؘ#FT���-�����G�ބ�6w8�6f�=QSΊ~$��
�Q��`	��n�7�o`���l�v��zS�.����ۈ���>3%$.�:�`g�KT�o-B�G���IrΓp�c>���HE�W�~ټk��I>��Gu�������,ZF1_��sB_��2���ٳ��N �Oga�q�?l�-hE�gq�&� �Xh�S,�L	#5���U�$V)ldm$���*\�_��J��� T]�Eqв�w���BMF�Ð��ӣ�t�פ�[�!���٪��1�8w�7���`�hb?�p���gl�W��Q�������U8�ۖ�ڎ�x����R.�u7���V����1N7d�J����Ԩ��Sp�遜�q�	�&Þ�V峬kk{�ξ�:�د���v��ɅKbJ�[΁g� �4�v�;��[��ш���tέS�s�b6Q����� ?Ȣ�D�wS,wOΖ�4u�Mt/�57��kFҫ���
L�v��"��O7�%J(�d� �Gg�f���uZ���9�0P|K\E��˧1W���*늒̳����k����oT8��v�)p0�ɏ]	rV=,T*�FC�%;����zd�
�O�wa��t$4��b]m�J�˕.# ��}���(�r���G������bb�;2Д�<Z [vte����Tׇ���T�����u'��]7
��	����c@�(��M�ӥ�x�a�ʥhG�|���,������Yȳo�5L٘M���p3ޫ�٢�&$�l2A��������%d�ۺ.���$z�]0'P3��7�r�:��O>�XX2;q����@ݑ�eɜ$�
W��^KO�@����w�ض��an��<?�9����e;*̖�ہ�F2@o_�>�%k����va?�+���y�Y��7�LƷ��M�v�$xJԚZ	 ����������B�h�ٌ�)�@��O5���fz:u���ۻ�����鷭ajM��:臃���!�,��ș�A�f������a���(�a٪L�C��͠}���:am�܂�8A�+{�tr����$����o��=B�{.
��q�F��1톘��_�N��)U��$��\+
W�1̓R���4`�i#4�9uo�;n��>#�m�X��ی���'>?;~	�n����'�u>1����UD�y�F�����I�$Y��"��G�EEL)5
p=׈!��L �O�����U	�VPtĞH�n����?G�M�"�q�;r���$}*d�!V@�S�H~ƥkg�ôF�jr,/͢���N^�E�	�����?�2I��i2{�E��U��,|�S,�S}���ښ\�ú��CF���^8C����9��O�:��ћ��G����e�a�d���;���Ԥ�O�W�Yʖ��=1�a�0֘x�^]��{P�p�t�M�Is|)/��@S.�.�0�h����~�\SMwC?E8N䪁4�2$H�C��غC\j��D���|����x~�:vj��s�"K��G1rh&$~�D���^�_k���0��Jq{����ZT�²��$l�.N��ڏ������U��^��YK2�O������,�U��7�S���H=m�~�pia��p,aR,�,���rܿ~����Wu3C����z�G�H�,�YQ�\�aCDR�T� � i�~���|�Tq�_�$%�"�g�/dD����2�d� ��At����P�,����'MW�e�HwYx�=�<7P��!���ѥ��
,Ӑm���RL��T,��R�!����4tN،?������=ܸI��8�-�P�<W��!�J\W�eGp\�r���Ɨ�~�,��bO�N׹P��c.I�?��9��/	�-5WCHOq��{k&Q��S˕ON�`Jo2��Ta&�N4_��sm�{#�����
)�o�;�l��Ol�;>�˴a&��s���4�2G�x\�5�2�n��隷�jI���3�J�H�r�e=f��:����M�y&�j�.����F8���������>�PX��:��]˪@�z�x  ���bL}׾�YJ�}��X���(Wj�:E�$����P�+�Ua&�>��Ȁw�A��"B� ?3�J���*�3��u;DtF���E:���sc��������-Rn?�A)��ӎ��xkO��Ej�\ ��P�5�K�%�l���51{Ir����?m��)m�NXȏ'��d���쯚0	�E��q�~d ��?��Bɋ��,�;���Ox)}�V^u�<�0ߩ���c�l6#p�9�ٸ����;:ټ�����k�q��1�'
�Ɉ�����0�d��7�띩p9_��H�|V_��m�A�zd<��*$�q�s���G�ϐa��w�1O��(�I��L���c�f�f��/{C�t��Q����q�_�.��%��A2#���=�@2T_ús�a`㵴͉w�K�����!�nE�G��-�׽���11�1z� `�BΚ�QQ�� ���8��9�Xs�*�_����{0o�GI����M����,��
(��8�C�n��y$V��Ք^̽ �͓�{	�)�_}�OZ������>ې�ꬢ]	��-��~|�3��,33��7��,}c�3�%��vg��2'f��B�/ȋ�?&~p#�F����C����J�Y�Y���z$�v�0�����.�*:���<�vl�����}�%���oΕ�ˎ�b[ƓS ��F�;��練n���	P+�g�i��k����W��J� ��lo@��@!Iы�bSG-.����|:��)}�0��:���c��p0p"��f�ɖ�٨�6J�cȭ��KCf9U.���Û.�L�K���cD��p���a)���t�T9FL=���{g�N�)H⦤� �����r,�ǔ�������G��X��k�N�ۓ/�ǬX&}���}a��I�i�W�-��_.^�0�^�~�rϻ�XrM(w=�W<6�j�a���J4@����3:l4�Ǫ�&z�mOc��77��?Ry`��B��`�
��{��WW@ԫ|��B���鞕���;/L�����D�$r������ag�n�g(�X��=�L�o?���nG���\�8��*+3!�SL���*��q0mVr�-ݛ���4�%�S��'F�gm����mr�U	>��ֹݮ$�G:�f����oțRZ��G\��bPX��&��}V��4a��8�/ի�8{�" �渱<����Q_�h��Ԭ��$#��g6P�U9,����N�H�0������ξ���"�z6�D�����7{D�B��?�*�����*��X��?| ��S!w�X��SOk\j�bфyۢ�<6����\NaF�Z�uԇ��%�ʊ�5�MD*��1(��t�kA^�Wjz���b qp���#�#���J��}+(߮�]@|����T��O)���ؾ��+r���Z1X��SJ��58���q����55bn�?:����f�;�#�H0s�5�Ց�k���Jr�꒩�x$�xp	�g�SZ#),�,�q=$�a;x��]:�ӧ�����%Ύ~�[�$ds�k�5�LD�f���	H���o.���!d2lq��s�뤞�`;ZzZ�'�5��_�u绲jV'l���FQ����'G�O��^T6�}K��u����/�X�������J�T�U�2(�8<@�J�kI.���d�����]�b�|z�J�0��ͣ�Dӆ���n�3~e�f̾�14><�P��W��0�f�g��cm
=�Ķ�?��)錐"��F���)�H��!e٠ޯ��n�߅%�O�β�!2�쁌A}I���kTG�V�[�UM�Vl�j:�������ĺ2�օ��}>�D�JϽ�_b'�*�����h��f�jX��.��ca�}�Ԗ����6r n"����Y�9�<d���EE=r>�_ٚ������Y�z;ǦP,r߱V��F�Y���v�)�$yv��w�l�w2�*]���Q�R`������]�a���;a��.��dw>Bh�?�5u\	��2�v]�<{�V�|s���X�1��>��7��Ī�zӞP��T�j�+��%X�����5Z�/?�I ����o���6X}�*͍���(&���X�H%M7{^��Y\�lإ��K�+?�s'@	-O�Zjq�P�����[��Z֠,n��������Xk�B�+����)J]@�w��|3��x��z��~�-}�Jd�>0o��K]OX�e�[d���	2.\�(��ҎiC���ki���x�Q�$��W�*��E�1�u��w����Ԡ|���KSk����PXZ�y����ۈS��W[��O�Y�:I�Bя�`��Po�k*�\/��Y&<l�G�u�~��쾔J �kܙ���=r��l�Oa��pnε�"�Ӻ]���y`-�G���`���PM�2HJ寗�F���G\#ӯN���)$�@�5��ܓ�n_���I�L�l����r���n}���}�J�<Pl�Zǐ�(E��z��O�JG'�P��i��'�\d�T���l���_z�t�n�H��󭑽4S���O����O��9=������/��/t;�#1UX�yt��x��!=�J)�f(�N��E��j!���A��%���"	���*ŕnm a�rM��>���o���!4��3�	,ùe��� �8�'NY�_i�WJ����ŋ��,�9�r-_�$S�*�֟g��>�u�g�o�3���ZnizY#��[��5��v�%ʡ(�A?���� taM���s{��L��8'��$�n���`TG������[�iN�_�q����>�cƖ��$���ZmZ����O��FA������ra��;�Ǩ�h���_F�B0�� ��F}�ȅ���r��M�OU����[;;כ[�3_�,��3 ��b��842��*�הϸ�T�0�rr�[��33�-�:��c:ü���)��e-V�9���rv"��q4&���BfT��l�Oj��/��7�c��GR�N��?a���L�2F������?VZ	��g"��-�O쉠���I$�y�_ʨIHw��;5���bH��
�oJ���	�Z�՟}(��Uj]��VU�1�|�A�"���u1��:s��
��s�Å�1%e?v0_�u2C�Ŕe�a�|g޵�V��\���6�O�����1J�(b�P<�s3x���g���x-a=��D��_t��`:��+榾c�aI�3١�����J�.�P���ډ�z(.��v�Ĝ�t�&�QBh�%k�tF_>���!�7�QVʾ���a��8��T(H���G~�:١]��0|{^�X��T��#\��}Y�y5[I���Le�Y&���k���Bd�� n�^Kɀ���W�&*("�}I(#׿�����9�+&��Gq)n�_o���k�����D�&闈΍ȨSC�P�d�w�vO.�Nz!hU]|g[ۿ-ٙ��̑�.h�����nD���mE��Y˚�]I�=$���X�eW��{����){�^�3�;�eּ���W�%P؝(��7��Q"��Oz��Tɏ� 6��E�Q>u봪���]5�糢���0	<$��RϦ�R����|�WI@��,�{���!���`M�y4C�Vy1���l �H�8<���[��E�����b��MD�y�6ޱ����[��s�%w��f�lw"�z�,����VhXS��pD5^�M:�1���>�gt����<�:9Z2)��� uG9�%�ۉh��e���9~���+o��qBM��'��ZyN�E�����Ѧ+��ӏ߹?%I��W
Ux`����,lD*��ZQ�E�4���۸�|r�+�mB��K��� &2����˾m�Y��k��C`b��̶�f���$e,���_�)
LR�w
����Fvs+s\8+7t:�����T�e�:y��)�X������l�Y�7X5b��i]wG>8!Z�&��5���%�3��"e�'ȩ�m~����7��i"l�;�a�YY�w�]�($��2\� ;��R��v�u����	Y�	���$�I&I�T��%��$���c�����Kb^%���]9uF�2�*mV����*u9 �����)�p�vзՃ�>��& 	�|��e�b���P|�� �5�o��/�*��>�~Y�1��$�����7����s�{��7�h�]���(IL��~ �_[�p��3WN�
��KۭiJ�C$�et���1%���t�M�o��p+�X{���^m�mc�6���e�Uv�+kO�sU�0��R�r`lTd�^�;v�Q�8z���{�%�\R����M�������=��)`+E���O���X���tVw|��\�c��ĴƨTc�Y��/�K'��YK�:/`],+(�
s����ܹ��_X�a��x��W�vZ�WG��2��36�z�T���Ԧ(�e�'��̐�d�0�
��Q�~�_G/���М���4to�7l��wAr@��_����g��?�V1�1W�hջ ��'���z�m��#��	B�@��9J�,!�z���U�V5�4�~*���;�T�Ps��K45�I]Pޥ�5����F�}h@'�q����vA�������b���x�;��`�d
y���+a^��W�ɉ���6u��ha+
�mX������IV-k=3R�˂�=����/���z`�)M	7��%^��)b>������ڍ�\5W�YԟnJG�2�
(�U�A�V8  �._^��%@K,}�q���d0@���	�j�R L� !�
%}vf�9�}잉�Zf�������8��(� �Q�b i?�e�Jb�l��::�M��ˡT�hx���m�Jȣ�Rf�ʭO��)���PLk0��,m}�{ˋ�}�a�z������#KΟ��D�l��p�4����0�)�%��{�P[��ԆM�@��R��dJ��ew�2͡�/�<�Mn�BB|b$,�ȵ�QHgP�l[	��ai�>���N�Ģ�5禇��4�^.q�uT�7ue���Zt�k�飄��YY@'�Y�~�{~�Y�k5k�Z���.�G�9)?�P�]ce~tc�vgV��W�v_/�m��͛��p��:}�|�J�WTN����!�W$* aG8>:5w:7���J�#����'�=��{Z��l�)~O� i��۴������7���(C_���%����+&G��{�#�t�ʠa�C����rraJHpg~��jOa�/+�_DOН$�u�q[)מ��J����Q�:����ZX>#�}����Y�A(ߒ��|��Q\
^Ygf�mmE���G���!���!�,��qV0��M�L�A�%�5�a���XKľ�1�Ol������Cfy�W�[{���ʼ��1y���Go$�01m.	l3��C�����[EtI;5�|r�d@r�����P���!m ��Lo%�YD�n7�R8ۼ����G�N�����hu�`���
,�W�A�ś��_��Ep�,<@eq���FG�s�r�R�ۉ�V��&N�Mz%U���"��Q��)%��W���WN�EU(3���I�/e^�&GWV�.����!0g��a��=a^T00����PoȺ��)��7٭S�Ș~;��}�l�'��I %e�rk!��qbv��Imx���`�>c�o#ot`rs�ƪǂ߲WN���fH�y�%s��k)!<���LU}u���F�%�N��Dw�Q�k@D�#W2 �M�YO.��Cw�t>ZNԚ|Y��}kt�?Z�N�Ό��0�>a�v_���̡�S.�̷Yf2t���=�nM�"�������,m�����CH�7D��N�����qT���i�K�vY�-����X�5Vg)��c@;����{!n��yē9��޳|�jl[�ܲ�MtR�8�P��%US��B��vI�����s���&u�{<	��]W�����[���>Jx��|*0&b"�����Iw��fz^� Uڲ���-�=�T$0��"S�ـD��z����D�]���-��F���i�'�WE��r�P��iJ���Z�7��ve@��&]8�ۈ����}���O���<��!˕�y�
����n�怸`q�^)�jlI��#ꚬ�	��j����ZWN��0��'��Nh�'��cZ\"���J�ͨt����똴~c�F��K�3Q��/�Ht�<�Å���*@��XV��w��1�R��C�F�U�b��ݏCV֤�ͤ2�N,l�oD��N�����㸴���Ag�Z�z�պި`��o�@`J�t�
�ʠ������Hw���������߰GfC�M��� ���~�W}daU�g�#���Ix�;��bR�7�m	 ��ӻ��9��|O��9~�'��*����䷏�S�
A!f��2OJ>r��W�{�卒��Q�n�N�(NI�6mD���o��[@q��QN�3���Mb^C��G~��3��
�,�o�nB��~6G9h�w��t�m6�>��:MNn�����L!ɢ>�g��#�Gٹ���t :��nO$1Q[���8���*��dbW�Ca�4�c��S�����NLbԵF�/��]$�|���_ �� sJ���-���	�y��f��i��^p�-K�n���:-��1UU2Z}m�|�y�m��"��H�a�#53��z�`q��2���īĄԮ��}
0�^]�����[,{]d,G���O��g}v�!z�t,�?���U��,�c�;	&k�g5ܬ�D�@�ݟ��pFzX��	���t����A>�8d⎴)��l��n: ��U�/����$��a��y�k��w�⊒���FW��.�C�s��tI�瑢��� Cj�IK�K�;g]}5�R6o6��`Dg��K�!oL��ƄO���4��~��X�H�q0�P����ϔ�{�rK���|O�O�m1�@���7��)����6fC�~���ד��A����ݭt��ڍ�����vc	��}���"�P�ij�3w���Y}̐���(�y7���}���@2:?:HE�)jG*u/�x����J���X�73����`܌2�&7�\Dٲ�	��64�fy�!�XB��	d�[\G�?�D����ԍ�i�3�����k��x�*��$)�52������d��o=Y�5~s:���َ��y�Y���S�"��":!�F�8�5c\��pvꘘ�p��O/���Hg��(~��5
���n-�#LT��+j��n8�oOu2e�J��)�Bd����M1�ޱ�Iw�Yn/�y��[W��Q�~Г���{�4��	�ﱴ���M�#��ʐ
U�Oy@�����d��.�!{d^�ũe�Ɗ5bgd�Gy��}=z��{n����9"N���t��L	�����S�99�hT���JX�L�{h��Z�}�G�= �s�J��TG���>|��WU�Y����1֨Vݱf�Q���3U%���M�?+���i����:��$�!c��|xz���m��N
�i'o���pPe�H��F�<�+m.�R�,�׭}�F�W2\֑���\e��Եr5]�螛��o���I�P�����K�i����ӡ�ܚ���*䙬���gZG�m�d��ZD�~�x��f��g���8�Աޕ��y�e��4��)m�g	���"�� ~��j��)G��nU8�qV�X�px���-a�f����P,L�v=s��<$��s��,Zk�&S䋫'4�B��H e܏��a|$G���9v]*�k�����҇���|�%M��}��=~��{���(� 4hz��e�I���:�{�ʚ>.���N�;�JU �C��;&��1����3dC�i�舏��,��ֈ�?V �(��z�֣�P��.��k ~Ņ<���X�D�G`8��V{����{%{0|�͵�e��#&/�Y3����/���X�y�۽z�W0i�Z��Cs�!���������R�@l�G�_�>�������I��W��ahJf�
��U`�b)�c̶(�6ή�:=��H5߾��c��dR���(7�����p�Q�եT�#C���J2G7�CD�h�}Д��b�zΥ���T�P��b��a�W�+9-�|���l���ͺ�m��D'����֤��5l�^��Ýt�:���р,A�ED�}af�������f��@�N�c�mC�P�@&A�)�����K����m���Щi]��n"T�q<�$2q{��D��ǺpZ#��	��/�>*~�vb����-\:]m!�����7�&��PS�������1$(��k~�����{f���5���D��]F����e�:�B���W4I}���1ʦ�͍S�m[�K��?fc�U�
��ȣ �u�X�mITyc��&���}>�H��N�,e��7�_����6zP�*�%����x�f��U.����U��j�M�Z����.V�kl-*�ow�+�hW��(X;AR��+�ʇ�Q3�Zo�����]�0�8���9����c�:��zYhZV�Fv@l��U�!P1S/�й+ҙ��������Cc�L�2���H J���05ܯAmiA�x8��*ȝ�FD\Y[nT���.�e��r���ϓδ�
��eg���q��H�!J��k��"8*��Q��z��4�/���Nݩ��\��uW�u1�H���Y�^����l�ّT�?�y���)���o^
�Bz�D_
��x�y�xܗO6��s���Y��j�|�q�W�.s�2��XK�|����+T���>� �Z�3E7ss��ag�e��4_���m�_�!,�V���)�<m��kRir*S�"w��8��� $y����v�eT�O�({PkB���
�n��/#�cs��?]~�r�!�Y��0:��a<�U%i6&>Swo��o}����:���tKj���ok�V�y�5�g��l�&��n���Ɋf?sd��%7Bl<�_ɫ����:�m�0��F�M��&9�q��t0�vΩ�8�4�Z����0�q(�����|���M��D�J8���o��ȑ{�~C�"ծ�O��y1�eJ�ϏH�� 2ȡ��M�c��U�@�]�#�j�~E�ۚ&c�T}@�H�hzm�o��5��#9��)����`�[�p��˃�)�˜���v�,�i7*D���_�馲���6R��ҏ�����y�����egm3o��D!���f�uͥ�=�W��*����%�dz.�+���t�ӰI�������(L>?{��7���SD
����Y����/���)%��΄�K�_2��X]b��3L��\*	#��D��˲��3YZ�,ﲛ%'\�vx�L��9	�JIM/**�Ϥm����WX(3�(�7���Q��Z^Q�8����N{b����_��b�of��buT�✈�8�x{��h��ʆ2$|:&�(���/��*��{��һ��)˅$��A�)?�ˌ�}�P;ϵW�	i�z�?��:��&Rn97�@v{:��maP�C�"~��F-���VA|,B4�E���v��tM<�N��e������7욇����<�4�,p�F�������4���+��h�i7ˢ��Hf2�<$�Ou��tW`p:�At��Au��L̩r�_��O��Ke�_�((�o��3�5�{��|��e��q�
�(�Zz�PZ<���B�{����B�^�fY�o�� ���N���VXd�9�ؖ�����q����]s�ܘ(:� �2@�����w<⼴AKط�|2���K���(��%4e�8{�����K%���}�r�wXY����8.'�-�;���� Ϝo�#4���+p���VdL��8�FvB`��U[%#輛$%�};v��L�
~�$��F�{�Q���^�C��r�w�)�C8�;�K�<|,}���N�Cj�M��yh�,-8q��Oh���%�	��׺�y�k�J�93�}�v����˶��i�w���Z�x����<s�1�m�Zf��V`K�~<{�ᢄ-��.Oi�9<2g;��kG�´�Un�.�#g�Gt��HxcJ���3��9^��z3;�v�喫�le]r	;���3)����\���i��/���u8M�@�#�@�͟#hk�E񭎕���\0+48���o9�s鏯�$�b=|״��CG�6?r��	���"DP�c��X��v;]�r_<X�xT�������������Hʼ�)UT��_In;X�:���0��Wq)Q��� �z�n�;�xf�>��IP~h}��~�,0I�@4�Eh��.t��`٢�Wm�i� �ːQ��C�?�M<�0s�#��=ŕ����� l��dL���˃�UV.�~x؃� �'oJ�k,���f�a��<�1Q�H_��!�V1ѝ)2���IP����W�f׳ȕ*c�ݟ�j�����g����R�L�<�~�h�����ctE�c3����(#�Jd��N`�t��0{����� l�+�����ڥ�"|eq4�����ݠbE����6[�=�)$��܏v;�`�'��|�%lCJj��uͯ"I�.��f�_��hL�
��a���<�w�½�[&�Lآ��d�-���c+du)�� �X@uP��i�D($7Y^���a;��V���;?�E�d7��*��Lvm�<��)" ��G�3^gP��f�ɧ�o���N޲�����P!�dI���h��<O�n��R���X��#*�i-Z~�Q{���F���<���!9F�*�>���Ң�!w�B���!5���!�Z�����{����q8���fy�u�&6��!*Ո���OM�.����>�h
Q�~�7]���ב9�L.�	Q[�;Ø��9�$���5�K�O��(K!��<��ۨ�ZLr,H�]�Ԥ�%zc�����E�Vd����b��{�����'���#-��<t�W�'��&\�UAţ��FqB 3a�9��r����0�s3]�*o�߾�ǝ˳�z���
e=�^�m�U�Ѫ|P��5���x� �g��+1�Ԗ}Ҽ�ߎ0��>�LO�F�����ýR�`D�Et�H{]�N^��Z����҃k�`�2��j��j�vq]�s�E�T�=I~n%�*^ߒ��7t8� CR{��}ّ���86������>3�Sf_�������c��CY�K��2����ي��E�R� nWJ ���{���cy{���X��{�h�AX�q�zv6<10@_}Cm���)w�*�]���H�7Y�\�E��SB�,�B����RxP�^�E(tՂ�t��s��Ӧ�!j�yA�k[����F|��
�+sA���bnQ{�#.��N�� ����;+N�r��`��*���� ���c����c�艨����*gc���9���C�g���g'�١�}>��k��"7�Wݽ3D�H��ղ�����m@���_�w�<o}dg�l)�J@Ez��J��{dN�8�%������w����V��D0�ͱr��s�{I��}�^'PMۏ����4�.���B�_����'��p��#�OL�T܌�ū8��u�k~iԸ[��蕴;(�%�W,�(ŝ�C�|�
�?C�|�����AW@	�-���_����\֤ԍ���n�k��V���l����^D��F�`c����[
��� b����`^�WM# �%�6��U��d��p���w���:����X�L�:�*��k�A0��8���r'�|�'m����r�&��:u\�F����Qcn�9���/3K�����q��%�~]�e.Q���3��hK��وe�>�í5�����	>Xh�'|26!�ی����(;;���\8J�၈b�k|�k�iR� `���*�t�A)hp{�,73⑱�b�c(g&P������6]4M�JFL�����	�@T��]Nݸ�o�Dq|K�L���1���{��Ee#3�ɯ��Յ���^�(�=
�׏R��Ȼ�m�"�ಖ'�!3�_�o�pJ$�Rc	�娚Z�;�����p��B@��=#�F��U�w)�Ƌ�!�4�]=�Xɟ�|��%i�pLlD�й�DT�l��_�W�L��n�s��8Q$�F�a��۳��p2��IfaLݢz:'g�v)z�g�Ξ�i	�|!}��"��������I�����,I`\B0V1��*��'����Ɩ���g/ωi��Y|��ڊP����3G��E����*���6Qp]Nѕ���rS�a4蟥��ר4����� baf5�Z�ȳw;�*���4C�Lm�� �#��
��i,��*�B���>�֙2�ͅ��4k{M���޻��%�"����Q�>�Q+E�˯)�J�$��~ؒ(��X(��d�S7&D��s��#@�Bv"��ۨ�q� �ms��-��*Tz���X�=i~r��O�:�u72 h>��(�����&K�;�̈́z��6"ݔ�C��eI=E�{.�dP���X�:b��+j�Q猕}���X�f�x���(�����#� M~f4u��p���2������F�t���ZR�ȡ��c�%����Ӫ�&% :̈=�nn���= J�&�f��@Z��9���1{iȮ�|E�[�M�jt}�u�x�=h���{���`��贊�I�2�G}�
Ij��z��\�a%�d=X�nC��Y"J�^��Z�s�/��E1���jt��Շ�ʻ�������؀��}���԰�ѺK$��T���Z��9$ե+����~�`[�g&ߨ|��2�X	��4�u���"g\`5��Q�;�d���;��r&��~0�>��»-Z�T{�a~g���a��  '��h�[�����}$�E��7:u�?b����Fġ����
�~��=^������6���o�Աk٢�|��LJm�.2�m��<f�R��nl���Iy�B�e#T8J�㯢]M�К�s��:R^�X~�O�K`|��G�<�q ��=���	�At���g=��jdy����6ީƝ>������=�ݣ4�s��Y5&b!lk��2��?G�Cs\DY�zZ�\kx�pg
��x&��"�;]��im}p�e������-5?c:L�?Di]j��!�N��ګY.+m�3��7r�7�LГ�X���<Q򑘨~����C����0E#y�Li �>�y���:�yp:bl��"�O��H�y��H%_n DA@�+�|Y����L/V
Ls˟ �W���s0��s�"N�<���Fw��`�b` �'��:�!B���w���.��jg-�_r��2*��(�2^$]2`�"YE�^�M�Hh6�ɗxJ ���jzT>���]�wƽ� ��'���x-��{��S��n\�H~��.�,]؉�*����X�8�ZI��l�F��N�~l��`k�ysp�X��ݑ�&��.H�ő&2�<��݅4q06���*��S�Uͮ����UE�}��seR��9_ֆ�=Q4"���5��@��(�[��I���ͣ�N�c�zî�0�Ӗ�
��\�R6 �P# ߸����C?p
�n8��g�q}U�(�����Af��hs�q��Qstg@�p�'`�S�F9T�#ސ:���([���o^[M�d�x����|n�f�U>��I��.�����IEtW�^��n{p^��nl�xP��`
<¤'����^�n�U�������M�F啅����g��$ʟ2��)�֢�4��|7��S=�g��w�T����Lp:f�B�;�y=�a�I���Y�m��A��iӕmuګ�!+��=���Ǝ��Ṟ��k��5D�`�l$c�6�9c����
��{oƋT{���h�u�S;��M"�IR�ϑf?n�ԽYo�V����Vt|){x�)�Rx� �;1�m�E:��g�ntb�sa�\m��'J�#�Ϳl�7�,�����J
E�Jt���r=��I�H"(��?6�����-��f����7NmdF������4����ޛ�x����|Y*� �jݥ�]0���0�Q�3�MZ���YP�3�௟��w��:%=����D��E�,ʨI.����)Z	{�����9���:A�6�~��y�@o�ٸV3ߑ���:+{�o
3�fy��^t7�^�O��L���G��$��	^Q肕6>n8�n��ke��Rmk8f �N�ʋ)�ȗ�^A�Z��)���L>ׄ�,��i�` ��S4�V5F��l����_���z���b|X���y�9��xJ'I��Z�2?:S��ۚ�J��@-��΃�O���{�A�SoE�}��J?5���))2Q��<��'�vK�����@�ƌgZ�z�FQ����p^�:'��{���!᱖�bb¹�W�$Cى������Ԭ`�:]�EA�a���!2��3e.î�Q�fz��Z��p��4T= ����oV/S�h�Y��"zw�\8�A��>31-[I��i����q`̄�"���4�]�P�(��S"��@Gˈx�>��5w��?�7�q2x�M�����3��Q��ah�D��ԭ^r}'斎^�3��"¶~�=gԲ�_1�`����yV=a���-_(P��T��'m���{M��<���U�sB�����BFm�8��b�&aA7� H1��гW%�L葇�Ua��A1q�L�]D���\�ZS�WG��"B`�|�lIJ���U�w3T|�r���o��-+#���H�r���ɒ �D�cDFQ��o��
, �d���+�x���̽�����{�Eʕ�g�{t͐��v��更�R��I'(�B,(�pa���X�������'@#oп�6@��P�>%��Rsm,x%2QXG�DZ�>�Ԫ�̽S��R�bwާ��Ig�;N?hf���*����
�ѷ����}�,Xٜ�]�R/7�rT~��0`~c�鍷�ɗ��cPl�gГ�vG�j{��:.�f}���1,F�־	���>	4��)A6���-F�����������py�QL�����<�G�} �bȤ�� H�E�O:��� 䊠|��oN����=\��Ml��EB��g�SM:Ĉ2�\�`��
-H ��%�k
���&�q��D1z8@�I�r%�����>�t>h	l��6��rtļ��\��o����v���ӓE�3:���Z?�^�VE|���Hpf���^���x����	whnۄ��r�9��f�����hS�Á �nI��ɿ8�O���7�p\:��}��~JRܠ AX���f�LT_��Ʃ�����6�B6Q��vw'�@v6s�C���ɇ%�Z\��ku1c�Sf
[o��'z���S���w����2�,�G`u`���e8^#���
}y#�g��hĚ�F�W����Z}SS�0Se�<eܞy���lI��O$C��۳�D;�P���r>�qM�w��f��@]��}�͇m��f=&��yOc�����_�y��?YW�1a�F:��η����8���x�6؈�1l��W�o�ju�q8ڐ�UN��������I��Tx����OyYD�l�A��RgGt"�]*yb;���oʡ����j����ހ�<Q���߈���:;�\�5�{�\�������/�'��	SP$��G�=�[�S�/�٪�ݰ�^*L0�I���t�L.��Ǘη4���i;@J=iKVD�Ȩ�Gu=��V3w+�d�;�uIq=���k,B�����:�u3�٨�e,�aoI��?�lkZO�^�ӰWRa(�q$���Y����$#D��z����fJe�F��K��%�V>X���|b0�ٺ�
q�宴�}��!�z'X��3�?D�����b�N�6��o����b��`��wY}�C*�������o!��*��{ow�T�<"�!vi�zW1����������OU���^+�y���ȬvI1�;y�~���4V�ݬ�
�z����1�]��hӭ[O_�L�e�V�D�7-w5?��ˮ\)�n1���]���� �(o@~]�d���Jac������
�YU��R`$�΅�]�#�Y]�Y�e�z��B���y���X��p��}k��|�J��ޙ�+>>�$e�y�����x�:`�~�r��������l�0QƧc'�0��PIs���$|��h�Xt*��c�@_�3��M�����N���Q8L
h��Ϟ$�j�&M�5=Sx�3�1ˤa����>���f��/��[7 �rаcY|�R�;��iD��;R4ʽ�H���c��Ç�M(Y[���mv��g��L��� ��`�9Ą����s�1��Ԅ�\zH��C\ �L���r�H�JC�74vc����q�I������O� n�C��e���C�x��gĘW�*�6q�����5:#�s��1m��[)�����8T{Ēcr9,?&ı`��_��y,^&�.J�e��m��9���@�m|�H�v�`T	�Nཿk>�pCl>�Tʵ@�.�f��ӎ������WZ d[l=4/���殄el�o�OgN2��4�0O��F��QC�<��V϶V�[����(?���F�<�Y��#m0�jQ�:>��J���
���� 8I>׋ԇ8��@fK���:�K0�4i�5���	2ތB��,�R�Ɋ.�3�}�[5 ��?�0�hzd��؉B�^�c�z���aWReBʚ
H3�*�&-z(~��,/<�����Qi�Lf�w�@�94,���3U.q��@ZC�IJLT�&G1�@�H3{n���_Jq[@�K�S�����"��~ȉ�K1Y���(vG-2��Djã7��s¿�=�qk�z�Vˊ�� r4��K����o~<��~���Yp���+i�zc�֧Mp�����kDe�K��R��h�
�>7���|A��e�<�bq�Q��\��#x���B� � 1���Q�6w\��ߙ���,�����}_�͖e��b����ݑ�@˶�!��%�LI;�|{d`�ጞ�i)k���=��¬�8R�M����i�3�Q	�-/�\��I��c3�� �!��rJ^�H0
��	߽b�(��Y�PyY�@$F�j�CZ��]u�R�ZT9�s0���<X�N�K����>�7�1��_�P��C>�+J�pz���ǟW.��8�0�8�]�J����΍�g2�O��s�%nH��?B�
C���\PSГ��A�h��0	�*��Q���9��pP��������gbi����tMØ�P����)GM�3~~U��#]�xFm�Xфe ���cQ6/Y�ݮ 3H���Eq4ahJ�g�-|�S�F�ҙ�U,��c��w �IV�BւF�B�4Hs�\Ķ|9��'��
N�Z�U��c���c[��b�V�gX���p�'M���u~� �C���A8)D����0��c���/lٱ^��m!Sμ���r�`�zR�1�!w!������|���V�S�,� @��gK*o��6f���݋�Vf�8��M����u��p��8B�������d���Ǒh^$�"��@kQD\�,��,E��W|�$2]�����g��︢�����������"mK��%V^T�H^�%M9d_e�~~Ms�����b��e��	�g61WD̒�z�1���"���ʓ3�f���(�.Ȩ䰮��K+>��,�B�}_�M��M�y]G����˚]Li���]�-�|�t�ם��GR�h�����ڐ+ԯn�H.7#�"�4�7_3b���/���_BS)� ��uEJLi�E������w_�8�hQ�7�����)Y\p���G�`���ѡ]+Tq�Q�u��oڠeru9_s��k���׃����W�NY��3^(��q���*�H���_�dQ�X�6�/"��z��P��� �ad~T2f���C��f��@ﵕ��pAn��C���Mi��,`@h��-
�jc�*�lk�սebZx�Ar�|q��N9d�d���F�p��?�����2�����6��E��os���w*{[�;��l#�iT�6��7~��_��=Ѽ�@XXrSoM�j.�ߩ��\�u˞����Y��<��r_D�������{}�����°s���f���R�;���q��?b�P�;I�<�)=�?�Ǎ��Ivלf��CQ��ƝE���|b�Q�sO�y].e}?�r��"��V�i�:1�����`���z�
�)�l��Ό"���h}�I֗?��N��L���B�'��0���Z�>gӥ.��ھc�������������ЬG���Y�G��mQ@�(6��g"ͶJ�:r�&��F���(�M��"�x�^�V�:����={w��[6Fn��MUr-z�ɀ5{���I8���{X�B�뭹�d/x�eE}(w�+�ը�������"GA��Ʊ���0�}��u9���� y����GG��%�g��b���N1���}�_�-a<���`�)`�'uR���ͅ���1���%hS�C�z��5�ջ,�DE�o�JI=�<<�A
�9��g��}���?�[�����t�[�0:�_Ɍ_�e��r����0�ɟ����
�G����#$��?�	���H�J-��9åY�=�i�2��j��%?��	��ɔOa�:MÝ]�F3�� �U��F��5�t������2'��X�_�L���k+7WG�`�Lq��En�1��s��P	��S��f��1���*���-r(_)P8�ks��<J���y ߋ������p_�/��^�-��	P'`Mፚ�{��8�4�܊�;8������TO}gN*���ƪХ�F�Pd�M���5p(�;\ݶ�J!	y�|���z�$�p���� Kb���<�R9����HV���h��D��]@�l�>�K��,��z����M�%��'�����ri@+�p�˭*5���|�q(�Z�J�+^���s�&�Npk�"�8tDk�-˰(n��F����L��i���@�O��z��{2�+RУ�Ryg|	
��7�T�CoW�zC˭�4$`�a^?d~uv{��;WeQv@�;k�0�H�	���o7ؗ���ϴP�$qq�˓њ�½�B؃{��]i�@�F��L�}��\ c�Y�B��4�S6���-���\����sV#�,���8_�<1O����Z��#9�H0�ѧ~Klǜy "� �5`3ck� �y�����/	dߏ��nھl|t#��ڒ�¥٪�����9���?���U��E��G�153USmQ�S��3�c�w����(�o��ѭ$���igB�e��iH.����i&��	��|R�4&���cm�%J�QgNe����d�i���M�B�%���ʐ%Y����E3:Z��m����L�ipp+�	XQ�C�
~n�)6O�X۴�ߠ�6e�iI����w	)�lQS��9�;���"�hY&_�Vr��WQ�c�H��%�+5�(�����v����ft��D������{.o�#���;	�8�
H�TZ�C���Q��G�	��&^M &N|�J��*y��t2�p�ql{zYP�O��~�������V?����L��Q�����2�+�|G��h��n<9շ~���d�Odg�e��y��R=s���`<A_B�E}�)N".T$�jQ��7�.��������Y�B���z�1�:��S�RUY\3��X��E&6�Y�E�A/�±7��!�6'�J~G~'�ZV��3ڒ��(H�-E lh� ���t_th/u�uݢ��@�% .����6�B�SO��t��XUJQ�[�G�@��)zަ\K@�h8�9HBMf�f�AA��5��o:p�"qj����\*u'�h7R/��C�([�a�ik������l|MjHpy�°
����V[�;7�9pܠ{xc4F����&)�ֈ���Zh��_5>t�s��ߴ���?��Hc##���C��_բ��l�y^��oT��F5�h(ъ 3 6@�ԭ��}h�~�US�kT��w�{l��
�t>���8j�Xe҉0.�� �Zfa��S.������DB���� <r9��pp�I���(�㤓�I*g��#��C� �}�Μ�ˋ��N�Ky��]Lv���P�z��P�2��O:�S���8~��(�rͲ1�T�f�bc5�b��Lљ�חK����S��/\8?qbk6"g��t��r�\���@w��f�`���Q�(�F�������1lO�L&��3��8ol��=<�@���dJ���d����
�
3�l\۸0:'�J :�~������.�.��iH�&N@L}����:�n*�L }�n���p����]S�2���mVG���]~.v�ry��'z چs���_¸ܥ$]�!E�$�8��"�>�@��o2R�����e���8wQ��Q8��X6�ۃ8�Oe�SZ,Ǯ����ǫ�f_�VSO�~�iIc?��$�,�Z�V���ܛ\ڮ;�U$�ŵ�� 7IvQ��ޚ���&�������	'p�^�wZWm��iVA=�&K��7:�[���IG��Ju�t�#����7�)��a/{l�0�v�9І�@���G/�aLS� 4[�|����Lo|q��~��������o+���q�Q���_O�F=}\�]�A��H����T��}y��èErri72���J��Ƽ� 鎍9��)N��d/�+�4�,K���ܓ�Z�Rha6$<�4=e|����Ym�]��o�~��~��-�G��~ 6fy���pb�{�Ƣ��i��NO�*���&�h͝dJ�S�#��u�H7);it.�2��f|����=ɏ3�w.i����횸�ܯ�a5���v��^�Y�+�qvM,�튡â��,�/�Sq�Y*
���%���N��ru"#��do!V��ɱ��fvÓhTMN(A���Ů�Hqߣ���;�0l(��1�M4\�PB���y�cy��9g���5b60ƅ�2�ݑW�f��Oac-��@q1{YM�������46tM�|}��D��7@E3E&��gj�=��i������ׅM	�
�<���%|���M֣�,HFz+ �ܖv R������m8�-W�>(�@���Q����u��6�ۦ�������÷)��W�$No��OY(��r�4}�u�8K(#�*�����dDT ���_�V7Y�����+گ�4=(�~�U�?K���``2A�f,UY��5n�ؽ�����R��,Z�d洼d��@�^&��"�H$	ͳ6ݧ���"���^�=$�����&� ���>�z����Ə�E�L��[sT �ʖY�y�
�`|��l��-��U��ã��k�Xc;[�'�6��l\T�_=��P�HO�@�dev2������$������Ҥ�0�5�ٺ�X�'�_���%8G>��\BYBQ��9����6�� ;ÇP#N�D5�����H���j������@orr��n���IAP-��f�"2aTV���;�6�{_�e��bE"�_1�-:��r�w7s��
�����ߺ�E9�x,?�^��껼��
��������s�0@u��4#*%�t ب�d���P�{O����K����[�,��?[�`��/�5=$;6��ar��~�@���k�.��P��15�O��T����k������UN�r�����>I<2��>�	Yh�|�_��g����rb����s����������a��v��ܡ^�I�r�4Z��~F�/-Ø��K����f�n]%�m���V�B)��6��, �Ghf.�`!�f3�H�4�L�-b�:�2%�B}��@�}���J#�@_�
ȕ؞���)�$�;Rk:���9��«خf�*�I���� ͊L��[�9�,�L�Y�o�^6~��P�Z��
��c訅5���Z�B���H��T��|��QdXE�΁�{觖���=�����]����i��	/a�)C-=??�U��{o֋�F������zLYg2���NI=oe���)���q�=�cڻ=�/e,�[�d�|���"����~�oe��8�{�<a/8<��7��[i�r1��'�	[V�S/�V��:�h�a���!Y��V�K� ��uϸ���I��.:�IF�H�Rr���x�Hz�.���p+��h��Ar2�
��SL�R�/S�$�e�!�sN��k�����X����5��0݌$������_hps�Er-)��5x"N��_{G��4]�6Ñ��9۰>�z�&lf5���$��#yZ��j�go��m��u�1�u;�����@3�\�����X�ɫ��g�s�o4�5Xit��qي{bÒր&0ԅ,D�h"d]�����T]KZG�j2.הu�D�`.�tud�����@g�F��D>��+�5@ى���m88\'
��
,�%Nbٛ,��N'���N>� ���b�/I1�3T�f�UN�!��e�b��׋V*Q4ƚ@5�*RD�v(D��VT��dڄ��S!ݑ��E�uJ��a��E�^�l�<���[0�ݚЅG�T�C8^Ox��g�_Ft'�;Fn�@�)Ơ(�d�үz���'����l�.q�Rݯ��˯)Ҝ �ŭ\Я}� ��,쮏���h����Ez�X=,���-�CnR�9�7��*���w?vྈRxvЀ2�O�}|3C�k ��E�H9�K���\����!W���zSHS�L�L5���X��/O��*�f��j�o���ܸ����4�j��\?���*��O�]m%�Q��xx��.x
a%	 �m �R����s�R2�B��u��86�Z���<��j�֛�n���d����A�'�`��58k���y�ԓ�zc^A�u��Z�o�v�yM��ȷ<�\���N�݊Hqqk�t1�VdцY1�[�����M�O��y͖>���>7�Q�	������Ҩ�ב�>��L�>f8�t}1T胸�z�+VK|�[űg)������+<N�F7����a�b�Hl�-Sqq����V�"�����U.�Lr�,�Le�䲎��Q���+��eep얄i;ey��H���Q���.�8�����qJ�y����XO�.�\�Mz,Q{i)����}� �N�쐹�03�X��}�1��*s����L���T#P�G�W�o���+:�[��t��C-T�bX�w<�(,������Ẅ����!S��JPu/�~i��w#���g�D�m(�x�=F���"rre|��_ɰ��w�^e�+Q�0�J�i��D�E�߭+�tp��c~�X�O�i�#�ԳJ�1<��C�Tb�ۍ _�����(�4���ނ�<���������D���Yyl��׎��_c��oQ�+�K���8�Y���'A�H:�����E�Pb���}�Ʃ��}u��gO����))�*4��>���+�=^�N^���-�g��3��`M�ج�i�U��:�/�Z?b����h)�@��GR�'��0�_mِY��qw��n���m t�����qZ	6�z.�����k+�b�M7�y*����I�����6P6�.��Q�^��Z�g�ʖG=Ӫi��c�vyu�,	�X9L�?hiv$ބ��!�耎`�X��A���g��#5gG��/ߣ� ���6�Y����ұ!=yb���M*1����P��,���ۯ���_�� 3V�E�D��;������G�/pap�TOZ�L��"�Xg
������I�h�=XU{XnB��d��\9R�M���;����w�߳C0:�x6%�������G��m�nQ�&�6{��P�~vkd�ő��������_5��p�07�{��U�����#��as=�;�)QJ���o���!)�f���3��ЕjX'�8���yT�r���H���Ji<?�(�lEe���q�8j���w*��\����1�
�%��9�4X�D���jQ�*r���x�iѧ<�d��b�^];�\T�彐,�(��y���k^�S(�k\S�y��3���9CVK'��IO����~K��d��f�S²[�0a� I9Ẋ���񎈒���x4��TZ�a��j7-z�o�a��k��1w�zd�q�6��x����D~��0�uU A`V#vE�s�.��^g2����0��ѭۇ݆OO���J�����L�o�1������x'e�rEi�*3�;4l4��������Y������:V��/�A'ۚdY���Nb7yǃ��zRn:Bt�ʫ'�K<?$�rNG7�ɻN�f���w�y��w�w��Ǟ>D�壡��:��[��d+a&��+�w韚j�#�<`K�k=����p�갶��;��-�e X,eʁ+Զ?�6ԇ����y��kW��L��1��k	�����ݖ`qNӮ� ��&�1ݿXw��Q ��������E�&JE��"{�ƀKr��=~���>Z�Մ��
I�8�����c4�󋪕��i�F�e��;�(>+��>�X�ӹ�CTO��tr��q�@�i�`����#Q.Dw��DLh���%�EG�ã��];���x�/N�P� �,I�c�ڙ<K�`���%m��w&������I	Η�G�Ռ�Oת�m�Ix�0��Y��z����Fe����]]n텱��2��H���62 s2�GM|�����V·��?a���uIǻ�@��@��b���OX]p{OA��]^VĒ�&�9��@I̟�֧�����3��`�6RfR˸��G�h�BkϿI��!�ǀ��d�'����zxt<Q��7@��|iw�VFy�ф=�N���=��4�v�MlI0c��9Q�s��_���E[���6(*��?i|}���D?�� �6�k�9Oou�P	�Y�!���w��@�2I�$�fN�~z^mj��b&�yx���Emڑy1�P7n[A'�}��h@S��I���h�dx�5�Lꄬ+��q�t��\]x�4|��:�gw�R��8 ��c�~�$#���3����\��֯3�;E���#�|$�wRN*��9h�7q#�4խ K3�'�蕪��N*�^[pn8
�$s���J^��.H��K*~H�K4P+iۆ�5(&^�o��8����W��:@i./�~��{I���=���YKa�3+��� �^���������+O�}�^���x�.��H]����q-�@e�����h���y]ǧz�pF��T؅�@o���!���2��2.jo�d���W����{��j�g��$,�B��B�B��P�#��NhԦiy�`a�*�&l׿��BJ?Iӈǚ�u |ϑ>w��2���ې�u�`~�V������pj��'%'���Wb��ٺ.J��2��H0�jG�����n݌y�����MA�/�0;�m?Ho�1��� ��C,�k�@�>F��j���j������M�%d���Z�xKCS��BÛp�S���`�r��r���gh�E_��j��b.ƨ�����Ѭ��D�w�E"b�/��o����^��TY���}��xP�=����F��Z�.X�Gl(i��R}�	t�w�Rl�eU����c��h?m�C�ނ '������'���
�v�͇6�1"�)�6��C�F,4+�|�l��D�ҥ���]on�[����㰯����/��&��%<�g'�F���&��g,�!E�g�,N��B��f5�M�x�Y�ht��ot�[�W_�hB6Ź��;<�<��i�Խ�Y��>�5���S!?ϭ�����M���4YT�)�VX�IE�0��Q�_Ė_W ����d�מa�=rɔ�ʀO,����a���cr
?o�K\~f�9�l��?{��&�1i��E��ES��6]FG#�H�~�����*썆�&K�f�k
\���rq�����k3��͵5�ڵtx]�RH���N*TA����G�'Ǻ�c;G���	SK~���O ��._�!?��V�KK��F�7�)�WH�C��[H���e$T6.U,>���5H�˧���F�Yĭ8���b�M�f�ܢ��
ЇLr�{g�uN�t�v�th�1�=��?S<m����p
87բW�$�Z��A'�H�gU��{��<5|E��5�ᰆLۗ�A���k��F�-�9I����m��b&����l�y$F7�C�9~h�I��q"KT�2ʩ�<7�=����}����v�4J��V�mm�:U��k;���z�b[t����D'��gxC^��U�`��ܰBh�<ZVLy��ݸ�;�����	�k�黙���7�u��_k�vC�yeSe��CS���������,��v񑞕��P��ˈ>z���� ����w����n��I;B��=���Q<g��@r�t0G1���A�%���J
5�,;�;"�֌��+/��fL��$�@(��m"��I]Y��������8�7G5Ko�x-3YD�� JthB���P���\��qe$:�.=�b%�O�W�y�9/�^�`G��:�u�4`�ɻC����A����/��j خ4�kٝ�p#�}%�u;�v	�_ �M�t`����E�D6� N�H�o3i����8�a�[�S�	gĻ�h��.K���m����#
l��Z��U�YvP
�QTc(��M�G�3��z~�ZVv����?!�#�;4�	�w�ȃ�g�yܮ�IIZBQ>����t_(>�>��(���o�2�/�{����%�_����$$������9�(�dH.ؔRU	�0��f�����i[�F�5|�J��c�uoR��O����)�|R%=o_�aq6D��9���xʶ[/�9�mMU5QAͲHl�f���u��)XJ|�ŵ���2���{�_-Or�F��
{����Qt�`:��^��#7;	�H�iHV;C����<�T���۩Q���go�h��[�7��n"�h����E��$���Z؇�nO:A"~h:�R?�g}��|A�e Q"��[�7x��io�`U�����X�i7�Z���ֈ����5K��d�{��0�o[G;�.�J�|Wu��6M�$����m�㝾�í�I��<�0�d��r�Ͳě	�c� %Cr�^���Tƣ{��8Cb�?�y~a�%xQ>��N
�I*�i�g*a��`���b���d���S5�Q�5�e�l�]kF�M˚Hh���T��-
�:xB2�;!R�'�fW�#��%���ġ�/�|��7k	sipZC%����Q�̕��3��������k��q������h�Na���>��.����9QͰ��j ��J��fQG�U��*�X�k��f0�(
��u�%�$(VC$��lcd�9��R� ���?p�Ѳ�e����kvٷ�9Z��4�68�w�<�������ُX�2��;D.�w�t��5c(I�!��yZ���r@r�6-��K���lWx����;JMw�G�v�a���U�Ƹ����J�O�'"ĸ��#�^�]C�<g�o(�ҒI-P��)[ߪ`_�M�C-�V>�E���w���DQ_'�"��e�K�8<���ʇy�`[��_K�5�e���7���%R������ߓ��U��Ŧ���4�.�V���@=��j�t�5i{��}�V�R *���qss����O�����N�RU���M��"G��ip��C�2�g^��ruAǖ�a�j�27.��
Q��Bt��6GU���)�#��[�b��FT���Ļ���[�W��vN����2�>A��N�k�`ĳ�ը�@�WC(yy�����Jt���~�X�$�%���tK��|��b�.ڻ�zKVBW�Gv��I:���n�������Y�U���ۨ��#���Zc,�t� �kؿc�n�YO*�o�N�1�'�Σ�h�Ĝ�٠A�^�"[��n��o<|;RK�*̮,g�N�����y{��L�%K[(z� -��j��C�0O��c������#Za<\�q<v\���������*Ş��i]�[W��x��a�f{�*u.Z½X����p�8c����ay��!�nxaBB:�|Ó�`p4^/j�r�'Vm�S�zB&[^g�g7�,n.�ź�ѸD���]\��C��U�7���K�^���[����E��N���A	;��u���Y�k�eci�3�p����:�]����<�˱���9�r�xGs%��Ly�0��6}\�m�m�b��mվQ���\錩��z�� �__�����p����"S~����,�<+i R�o-^Q�ַy�'i�Z����hf"��pǛ�5ƈ$����r���ܹ�c���uq]?M�
��v�Y���"8�3��y`]rWbw�����d���V9	D<���b��JP[ �:��Oif�˗D�֙�V���3?mX��x�5���[W�������&�<����v��"!�q��$zd��jk�V���m�u/�װ���A�7d��D�����p�J��(d�lևX9d�q/�I��s�	4�j=��yڰwM'\寢JMk�m�����D�}sXXؓ�d1��,�^����y�v#nQ��x�)L����:�7�����ZSHp�Y0�b��f㑿�gqs�2�0�DJ��*[#���-�j�@���nv>�p�B|�BdgB�E������~�l.2T/	�1YX|���xU���H���95l�-���Z�=d,pk��^�Uwo�J9|S՟�9�z��_�~���]C ��L�O��R:<.6�~��嗡ai�w�5��ڹ9S�M.`�^L��mi[S������Ys�lyJ��݄�2՚�oi�J5�q�g�������п��;O7+B.����Q�|Լ��3��:֐�N{�ЎJXH�Rz���ҝ?D{�u��^4)9��"��`tXo����։��F�u�� �ҭdA�\����a�G��ȘX)�^�����4o��W�����`_H�j�P���'k�&�2Z���Y��M���U��R�)k"�T��.�{?�e�9*8d27�v~>���vH���2��|���Mc� ���ԄI��; ����y�U��7���=쒤m3�����o���2��q��a�iJGO�{`��݇��ș��1��୷v�+s�X��|)��
�L����.F����Ȯ��jg~�����<����̃�����<c�N����c͓���dH�H2�^p[޺�����C�t��d���q;q$��\7LO@*���u했�i��ҋ�N�����o: "���JrQ@�	�G�L5��p�\kj@�&ދ���g_�Xƿ>+��r%��f��_�5��_	I���� `n���^T��W_hHKc�NR��"���gq�~�{К�{�پ1I��9|a�<#�% ��OIAff�����i�SC��:���P�N��l^�:�&(n޿�緖�����H6ϠI/�dpa�e���b��K[�y���'��7�%o蛟�L��ܯ�_��?��D�%)��@�a�{�� �l��?��
�+M�����O�f�VB's�>�ܼ�����p��$�O���䬬{`	j+̶��XvS�EI"L9I%}%�;i.�lEی��bC�c���9�z��#�`��5���=h��22�w�ا|��?�a���kĦ$Yci�����[�m^t-n{�V*�r�F�7�F��d�_Q���ۊe�yX�˨�Q6U�7�G%*ai�M4��O�U�ߎ����6�	-"�H`ߚe� �FI?�Z�Ԟ�����S)ϙ��)���m��)�vh"D�/���*M}W�fN����b��]|��?y�5c)����y��J����v���5N=�3��`�G�a �]Q%������o��_�a��I!{�݊=���l�^Z�6��;���+��L���B�Z_*[zٜ�h8�q�"�2���
j��#ァI��1sIZ��#G%��`R��u��VU�-D/�����-8�n�� v��\V���Q7��K':��s�r��g���_&�JX��7T�$o���FٲP�JlG���u"�J*��l�A���%��o∩b�߷�k:d4�~h��}'�[e�2p�po�yZ"j�
'?���.�z8i���ܚ(�³3���
�uUO��1��g�X��X2�E!���uX�3��1s�`/-��ڒs�#U�K$C����f����C����1� �Q��X!b�ˋ������'��A5v�ޘ�j������E�%�=�������<��|���.NA\�WM���[�����#&3��%��遾�)V�Y!^�:�5�zC�5�]?��uт�ܑ���,Ȳ�i�����t�l��wD8��
��H�1OJ7��@E��%����,)=�����"	*����e�ӡݛ(dK�b����F�rkđF~q�1���
�W+���b��#U�!8a"Ar��4���R#7+�0:a5�.���ʀʚ���_��Ea�HHIz��u�t��_��[t[�)��+�� ycKF2Sc��*^��7ze��2�n!q���1�M��Z޻�"k}ㅦ����0*J��W\�����_?����ّb��E
�����H��D;j�3K{��&L�|hzF�M��g=f?����5e�?����4���sN����|M����1;x���HfK�ռa� H�,ɬ|*GL�H��� *3@:	�H�Q�SÆN��'C��;m�Y�bS�����d�w%��}�ʴ ?r�M����,��9��ፄ`��1�H�L�״-+fk�������A��xp^�E^I#�s���_$�Pa�qvF�Hv�L�7'��51d}���y�7(��tnJrc$�x�4��?�ߏTk�糥���8�eڙ5�M�Q��d��=����l�;ɒ	�[i��*��3ٗR(X9�je#��.�V�I��8N�a �����qI�ʩ	��ݻ�A�
��d�V>��^7Mý��"6	Key�M�i�4������!����%W��~;�ߙ�Z�!�a�p�t/A�*�:�.��"���H�<��d}�P$�e��6I�Q?�! �	c��l^@�2�+�H��Y�yQ�5���ė��rC_5�ؠ��/��ىќ��c��,�/���:˂][cZ"�C6d����[��9l��w�x�d_�gӁf`���K#�C��>T���Y"dz��͓��E��w�!�����}���%[�"�x���w�f�SsA���S���nIph���b����f�? 8�}��?��-E�tD��?0�6�����M��UGhr��v&`?�
Ua�����hRݬ$t
9KԀ���8[t�JBw��zQo+��-�y;9"����=����4����N�s% � �'f��Pw�{�0�8�f��~,,�:
ӏ�~c�
2$�i&���C� �zl�g"�X^QV;S���G��t�b7⢍�
8�B�������n�\� g��q������������)|U�e�������ph�\�1���ÜW�ME�+�vO?��O����IE�������(�^g5F���M#��c��CQ��OZh�_��ߌ!���S�l*}���;�c%�j��)9��ŕ}�&_l/��>�o�S���J�^��0�ℹ���ǚn��m~�j�=z��m�����*��S�ϱe���"F/�G3 ��L{�Ĕ�I��/[�������U����C�Ld���G�5�*��X�t	6�����;�����_�$����!��~�#�L�C-��ɤOz1b �ϑc��)
��^`�Y��H>~@�~�K^���ق����.�lf7�X4u�� ��������~�e�pg)��	Ѯ˺X�j�HS�����){#����8R�i�`N�	����	H�TmCX�x�)�2����'*����)|�����P��a>	�[*7�F�JTRn�*�L��'�=�Tq����	�������A�1!�Á�>�bÒJ�$��H��)�t�4̷���_��"!��0Sb����mԱ�\V�1�j�nkco�!J`8K8э2���,��~��B�w稱�SM�U��I����13�>#�_gZ����_�_�Cy1�B�y��9~h\��.����� e�X�Rt%�X/����7Ck�v=E��Ƃ=Y��u(����@� ���z�.	U�@BOư7G���\�����C���ѵ&ޢ���/>�������	����6���NيCG>�CDG����y�ԲΘ(��ud����G��,bA�~�T�?6�X�|��\�S�1SЦۭʺ-��!�D%��:����ra*�:l�������׌��T~��爵�©=@����"~��&�c��޶��H�7j��<�1%��O�P'��,��GI�NyM�X�9��V��.O�M�B&�<H��2�K�&�����h%�_�m�uSw6�5(���;l�;��C=�h�ͥ���y�����ņ;eN"�J��6���(v�|����p�۫��y?P�Q��b���l?����giX{Ou��lT�=D�^S���N���ْ��L�Ҕ��3IА���A�J	n�t��Z�|D;b� �qN�<L~�����bg�	��HK^���F)%N]��0����M���y*��}��l��=oZ�|��9�[6z����v�s��'��iVC�ӧ����-����)��sL!6اO@�U����,?��bp��-�x(�M���sr����&DڮW/�+��Z�ypf߃�j� ��k�'D0���[�����Bd&�:Vk�����ȇ���ج�P���6Q��"����G��5G4�O���o��r�D�%��:݀�b�?�d����&
�B�:\��\��u�c��ǹ��x}V�����c.�@�L��
��<߲� -��p�Ue��Is1��jo�}����b��T�Ì.WV�Yۊ|�"�4C#\��&�~�C.,b������4�x7G�Y-N ,	�g���j-��I@�tl6�<{5a���B���z�8��樕�<�H�~Y�G�*3Q�*��l�x|5��9�I"됖b�>7�ۺY3+`��UD��+-���1�`�㽽�X��5�p�{R1��O-�A�/�j1�ot�W+����9�d�D����͟�Z?�fLNQm�=s|V&�D����F#�C��B��"y*�f���o�|��^Ė@���	�"Q�N1Ɨe?L2T�meZ��5N��f�@I�p�$��|K��Yp���A��C�	n��:���=|�ʻ�%(O���~5�y׫�a/vyi9��G�*0��R�&�O6�SBgo����"�Uc�8ݞaY��	eŞ	Z�������TZ,	����E�lu}�jo��dW;�B�,T�}��CeWs��Fkܯ8��A̔x��Hi��9�s�Ԅ:��<�h��@��Xl�)�
޷9��LJ�u�c��#�y�D�)�w��_�v��c�ݱi��"섷¾fn�hw8�<�;�T���q�;�N֡�Ȱ�Yth�m<Ŧ[r��.X�W�\��d�˰(V!<mlb�P�w��<��EI
�?R������m�[�{if1�8m��n��Ʌ�64/���%Ԫ�ITٓ�4�6�����:�`&ԩy�PY�SҶ�r~���r��VZ����W���kH��XC�,����������~�]}��i���)(2�ΉY��;�N�XV��y�ݒ��M�v�.��a��a[� �?��L�h����I��)"(�v"Q�Ϡ�)��w����8��7�g��_ES��A���F���|�X�F�k������B��]M�x��	h�+�k��X�k�/Z��U�	.R�MsKǬ�R�{{����ų�ﳵI��n^�sfG�8�}��vOL�Z�z˵ �&�A��W2���	��`�d�$��Ǔr���|- ��4g��7��%*m�������C���CZ�b�
�V3�iv�4�'t_�/8�R�¤P�g�w!�0K�Mw�]"e!�B#��2!g|&�l<&h c������)S�F�3>4���a6���;�������i�0��e%�Q�F_}9ؖ?^@¬����ìe�MN�;�׶A��F���0��M��H﹦���u;�F�8���m&#��Sk��?��29F�ml'�����c-	&��4�v�w"���'�y�苶�lo��Yhڅr7�~䔖� ����^��/�{�ݻ��<�7�4)��=���u��8������̩u?amO�yn?z0� �w˝ңIC�c���z?nr�J���ht��c���#����b�����Kg�?��g��?8a1��I�� x�uSK��i�#y�+&�z���ŭR�N,�z��#���u۫�dsn�τ[�+@hr�� o������v6S�ԣ��fhtǭ.��D��1g�n��ϥ���δg��=��α`ԝ��U�S��p[響�.��|�6,ʖ��C�J��L5�͢q���m��򿫐ً8߷��D1��"�]�G��E�4��Q'�*�.�{�`Pw]�ت�raJD{��4y#�����px�l9�ep�:osK.(��2�P�v$GU�H^o�E-Q�.Ol��I�Kݫ~hGj�/�r�H�'>S�\9:%�\$��u[7��`kLI]�!Zn�6}��XZț��K�v��s��B�H�I���%1���I 'K����O�#h��!�˪�e���6�W_c�����b�u��[$x�Z��I�~�4��=?"�(�.�I�+��/�I��@��p���#��&lC�0U�+�h�a��4G����[B*��1�8���֢6	� Q��� �%�B6�� �-����E5��g�-�ԙ�T�3�����缢�xn���"S�s;�%0#ܟ��8X��m9c\�ZZ�M��c�Ab����EW��W��Z�k�OP.~�P���C57���4Tx����U5b��Ƭߟ� %j+⬶Ɋ7��o������OI���5CZ=	���`0V��L���5!\���/��"JD�Ɔ�z�'8�ݼ��W�^lv�gl���f@���]�ݫ���!���Y+.}	���6&��|�.�F���J��Zwh9(]zڼM�w������l�3������^4rﭫ< �ge�?oad��<�$�ԗKS���j�(�wYǓ��~;	
�����_�A9�J���ۘr���䠛h�Gэs���ҭ��&QR�Pa�]��ف��b��O}����!���^+]�!�-nJ���Ė-�_!��k�.����(tN��â�3�I:�=�^��W�o�%[�{|��X��z����a�{|��'eJ�X��1N�jl�p<�M򗬫*'�䣐l'��ϦmޞXuҹ����0Ā�J���+%�����̈&���2F����~i]Rl�p�M8�9z�f3rM�N�b&�.�,����'3m��Ĩ�hY�(�=����&sy���Y~U��G|7L{�3�Ilu9Sa�&�����#ٺ��(�<3I��!R�c-�����0���H��^N�Ԝ�\���a�RΊv�ه�_��VoJ�h<�^��X0���f��
�t'�ļ��x�IZi��5 |�.���PY��RD�n`9��=��e�`:Z���2��i��j�Z̳�*�_&�V��ۃz�:x�0�>���B�i�I��{�� Ot8�Ĭ���ߢk�6 s����qM�&�e��p�K�c�*�6h-���&�K��}��&kD/���O-��4�y2��똦��\���&:#Nd��^6�<�dzz��oH�X�m��&�fx�@l �BB���~�T��|j\Lk��$|D����PM.�o줿��Y�3�^4�# �4*i��Qĵ0�h����]+�\׸[�97njC��m�:���t���� �iY��cx#��i,���.�t2�l�� �;Z
3Y1���P�_���1��ǰ�ɤ	$�p�1�v�3�=g����Ύk�F�S1��L${.�NJ��"���g:�i����?󎔲3؂F�w�|�̫Wa�m+X1�0�:x������XX�߬漎���%$�}�~ý#�c�Y�D���Ȓ���u�m�B����h��af�]��9pB*��xf�u�����w�S͍���q�!T�\Cu�ӕ�8��t-�E���Z��&˅�`o��Y+��@�<�c����J���_b�k ��;�6X�~h�QvQҋ�G��?!�j=�`�X�`�/"��o�*R	q�����Z��l�C^�h��@��@�'�Ig,)"Z�vШkb�6R�s�����:�$��>�ҋ4�j0�)�t��a�yǖo�N������U��XIDJ&� e�@�#��|���������	�ǹj�¸�	�@W����L��'����q�����{ES'ΰ��4�d� ��&>I 5���<�Gh��s����cpA�U�����L#NM%r����h��ņA
/�.9۟���{�j���s�;�GJd�t_�vN��p�g����,�Ё���Q�P��Wb��SY�ͼ	�eZ�=�ר���U�Y��C���橷޽9�_�/K���%i�0y�:|�
��8�\�|K�it?��1�Ȑ��c�
(��[�V}�d��?�W���eiŶ4��)Ė�HX���3��n4���������I�'��͑"U�3�D���D�d��U��|k���]M�8����NZ��Z*�g{�C�L�[��1��M�ً�jFg@ xP5pr�A"��Z�1���7�� MHGU�ZY�3֡A̭�	W.�'�aT.#\.\3��y^`�[ܷ�����_k����z-�q���N�ʫ�2@p��cG�!����E���ׅ��v����_^�5/��W����HyT+s��Hz1��^l�˅�+���R�����j���^BT�jڎ��G��j��ł[O�h���;y=�v����v�6�R�I^���W�x���Q/�m?��� �<��#>�&�qٰ"w���,Z���#/媉\WW�D��+9,ze��� ��!��q'n����(�v���� j�T�Vpb9}�	�����
�ܔ�D5wN�%�~Mp"�H��|�a+��Lk�VS[Fڷj)ܣ�Ӧ�O���*�p1}���_����s��@'�]`a������ZBO��K#ϹO�7��c�}>���T��~7j�����jz��4LM�o�39���w�)��Hf�9���St0�,	���)C�a�ۖ��(��4H�j[��멓'nk�#홡h>���^.�F�MO+�;�No]k���ۅ��%�|̠��\H�`*C�9;Fn��y�~w�|��9��������f'Y�	,�>�Wu1N"0n0���5L�����6�t����^ҫ"������Q�5*�;���#6
]QAJ�
�s�8xx���W��v�w�BD�{1u%�D�}���8ӺY*<��F&���,�%���O	��ޢ�*M`-��I5�qP��(W=�^7j��\T'sw��#���=_Hc�x���E�,o�#vFpo[�ԙ����.��σ���$�m��/��Ɏ���A��ݎ�����΍�5�L�y3PkV��Xe���Id@�ꀡ��E���"�Gf�浩���Z��0�P,���,�g&�;�Y�ʽ! B=_��a�D6�R��`�n{bbȰwS�m�Ĩʾ�4Լ�(�%�a�|�֪�-}3Ox��miZ}�g<s��rl[xEҙ�m9�����m��v��p����0)?���[�0{ ���.Ƚ�F�{��M�ZGH_�hi:]g���8*s�
���|~j0/tB8j�փ��ԫ����	��w:p�_6���CZ.�E����ä��ȸ�[Z���'�)��7�xn?C��k5��]���Go������U�}���/�����P���a� @%���;;���
M
m�.?��lB��,��>�� P�:4���S�$��qs�tnzC�0Eb*���
j��"��ߝ�(�e��Y�S�T�6Rq�f�h��C�-!q�?Evp|�XW����<@� MP�"
3�Z%���+F��� ���]|eL�X�����g�KH3�i�O��W1�5�Z5���Ol�k`��lp��gP�~@�l�ʣo�F�.�Q�8�d���k����%B{�hu�^���w\D��kq JF�< DI�j���RS.�aG�87��t���&|[7�6&��0x�ۤ�75��u*1\&���;�)��a����D�16�� �a�$�f&�ȫV��
��v���9Ǖn;�!?������t��ӭ�l���ݬe�e������s��؊Yg�R.Ťu���i׋�|�,A�znebi󂳭�`y`
�B��޸s�m&��Dc]�|z�qW�>su��k:���Ј)SVYZ�V�w�EX�v��r�8�*�P�em-�Ny���sY�I�A����u���F�� ����`��9H%��pvs�oڀ��>g�/9�&�����E�%�H����k�_�y7wD��$�r�BH���Q���=<�cg��"�"{ېfMP�������`j���kW��hvt�� ��HTc!���Y��V�IX��Z#6<��a�ꡈ��k
;L��֛���0����W�U:�E�tsC����A<fN�4e���>	���L��o�A����}��~�X��9B6'J��_z��yZ�|r"�^toѶ����^&���
Y|���n��'�K/������ѣw(�|-�밺�,��G?�=���-It�19	�ڂ��%4[+oB+�y�t��	�H�&�`�������H$���Ѱ����zUt,$�0���F��)�J���4[��B���ypX��w9��B�lRV�j��sQ���ܼv_pf9� �Oh�P�Rz�H��o����⣃�3%�m ��Llɽ$�h`�s�ug�~�=�����bçO9Hy���ع�?fR��&/�H՞�Um�ТP�Y�p[��o�Ţ��6>�:��K}vt�'���Fq4��P'\t�*&H�x��p -�mOY,���s�=�	�6d��Ў7sB�f����G]fJ���sO�D�K{fa�883@?��3��r܅�u�x�r���$��l��m�����ܼ�i���Wۍa�<[d�70�����C�F/���.!F�AKCx�����l4v���"��+��r�cӻ���8�.�m����o8�e��  &T4����2VV�}��i;ݯkd]b(U㯭BW��b�a9�/�9r���ӏRVE;�{*N�]ׅ"�УO�9pIE�m��
~�R�!�.!j�� ��,�ְ9�z��"�����w���cb����?��? �a�X"r�nj
�X�]�*d=�%P�S;�n��6�}����fvQ#����>�z���������2��pGO��!q��$��$oJ�mgb��ʶ﫿2�3����@�jV@���+��Z���u�X������i����J��8�rẺ�����拏g,4 A�V��Z+|;U�_rX3zb��T"{?ȏ��4��o�Ѐv�
�X�|���1X>jƥ�Ő��o5c���{yn_ݾSL�X�̿qAO�d�`K�>m_�D���j��-�x�9�7��.��J������,�~�����>HsD��E1�f�P����k�!�h6�HVe���������_���DQ`fT��ջX��bO�Mr ")���[O���y|���K~�;VLVN�O��"�v��7�5��9$(�:��V�ֹ�o1Z���Bj��]�:�N������*�Q`��n&� {'���[�� V7�-�Y��fwN^7�4��e�l�>�ه���Ҥ������Q�]�����	ˑ�_=�_�ޭ�!�J�=��A�]A%�ئK�WE�J�l�?e�\al[�B�o�U� �Se��Mu�Ћx\\ة5�,l����.,m�ڐ��qo�y<��=!ϖ��G8�_�D������1�̫�U�[瑗m��{j�7�����^�/��M�-��VP�ё��cI�qk7���n�~�������MZU1�{{]3ß9]���_K��v�KوamgK��a���N��}J��&ɞ�ݷ]�t]����ǮU#o����� ᵱ��TD�^>�+g�)��U�����U	�����m���ۂ���*ʌt}�-A	�ItE� k�x�����WBθ}]?�i%ի�U�\ x�ٯ����������K��i������GY��p	�S�C�p��՘i0�\T����$f܎Ƞø��҂<�����8E�T��J8QC���P�5��;������X��̂~*��j�k0��\����[��KA,��G��e8�����"�pw{:ț���Ê���i�L!���I��?!�"�ƙ�b��{�F�m.�|�FK��G���ɦ�q�o�&��<��{O�,eM��HjH��AP�M$1��L��^9��}���T�\(=��o2��+-��E����G煀ƙ�"�,����F��CJ��А�4�2R`cG@ZN�68�6��xU��?�J�v�mҨ��SZO]Mz�a�,.�w���R4�&9�ށ�j5&�{j�}��/�/��F���N�Uױ.)Vȅ�f^z�Y~�����O��j)�d�'/$��P;��� (����_����MQ�?i#qZՔ"le��VI�$8�cD�o�"~�pa:��B'K2�2��R���O�=_kZ���`� ��J�jh3���x���e�!S��ݹPo)40f�ʈG|j�r��"JLv�s�r���eb�� +x�2]p���$	HE@��Z�M��\Mʨ�D!+
pT}��9|EJs�r�$�^�w4[��-bS��Q:��䣜E~<p�0�����0��;�}Ρf-���@]�J���¡q̶݊��f�pvi�y�h�r#�a�{`�b#����q_����򣮞�$�Qo�o�^�;�Ĕ��ǤIB�Ԁ~�X	�n2�\����/fl�����]�J�܁x�.%�)���$V<��x:Z7��pf�2�>%I?����I#])^�]I�>-�z0u�a�7�% 6Z�$�@7�2�,&B�~E�N�y�qՠ�7�g���V���i�c5KXk�y^��wۙ�ۣYcx\��V��F�J�F���s���2�fFo�SӚ{I�m�覄#%�5.:�Hс��ω���Vi|m�|��ﰐ��1�e)�9�n���M3I2�_���JL�$<�x� S��7��ip��lw����U�����h��4KE`#�HO����E9�}���Z���>ͫ��5Y-u�QH'׊x�6\}�_���4Ȧ3�2��p˜	bD�ķD��)��-ǈ�S��*�a��n�)�s�W{cD�E�уU�nO�H��N;�A8���"a��N�l>݈���~IU!?q�aa��u�Ȯ��P��o%wVſ����[�;�� ��f������E'��D��T�%(5�76������Y�8�1y���;�纂��Y�mb����j6BI�fr-=��1M��6�^�����:}�"��=�1���:�N	F��6�\����ιMYtu[M��Ȃ������U��^P�8���/a�B��A�h|��u�ȴ������!C�����`�X �r���l�;�%���)#.k�C�X*.+G�K��X�:��c�Ѫѕ�!�E�&	U	��%Tܚ	�OW��&���b+@�e�9��{�n�En�Ls�6 ����n1k|��ޮ�DB�xfn7�˿�X�xE�[��	���k�3�p�i��u�@��S n�Q�S��w�|�'gGo��� AO]2tx���2�y�^��󳺫��nv(F���!�kt׈z�oc��ᬻ�L�@ <�i"�啵b>Q\����U�Tp�����\+�A���w�-0� U�*�G�/��	�4.;�~41vPi�ϰ߅���j�9�͑3
��.�=�&nY����?Uҗ�}w��Y�ʙ
���ѴF$24����=<&���� ��m��gˁ��lx�?X<��	ewa�離ٌ�J�||���]�)��i$�,���dn�I����/鴜UUMp=F�Z��4��v�d�qoI�s�s��ʭ+
]5*8�DNG܂4�e��,�4��b�c���S|�$�gXH~��i�)�֨�Y�>C;������vKP~�yz	;s��O�D�꺔ix/�<�tu�@1{e�N���n�j?���@�5��FT��������j7T=�CV�Ri�t���Olv1�.��k�hĞ�'�p�]o�q�}T��,�rh�
�> �6�jm�z�R��+�{�����P��X�/�V��V e��[��S�P2����� 1uh�dX�(.n1{x�D���4��������z]3ߢX�g�ɰ����hE��q��#諩i����,uԗU;__lV
spr����b����ឮ�c��@'�a3�v�$M���!��yӺ�����i۩�����V���a{����S�~����"Aɖ{Z�:��NBM����-�@�A�
)	Y���#sf��'��0 Q�V&�I��*�^��JjG�-,�Dx�t3�}5r�B��C��G�[��_�|�rfJ0�٣�E�ɫ�-zZK*�^�+�ߵuCo� ƈ~1?9�pu#O��j����������sBv.4��J���ſ]�̎9y%��H���1]�I����ޚ�|�1SY83�ԣ� �]n$-�b����op��Oy�-T��Bn���#�������fT8��\�Y�~$ڭ3Ǆ�5:��a|�Ҵ���Q����^�54L�~�������$<D5�z"(���'���1�q��C���%��^�
��"���o���de䍾+���S$���0DO��m���p0
q��iy��ąX%o��3x�](�,*V_Z�*��~�5wٷS��=�rO!n� |�u9e�w6G=.t�0ȇ/�`@�Q���ABn���	�>��dJs�j\�7c6��"���g��m�`à~�ᬶ�巟�[Z�FN&{�
p	g��F��4��a/��A}���=.�7�Ok�N���� ���Y�?�.kᙦ5s���#�[����u��l�<�0�8�O�~3�&����R�����W1������z�p�9L��W�*��`p�_�����L9a�ָ6sCj�D��)���O���GX�SWK��_�l�L}Cf-����<�h���rF�E��-]�.�m<�������c|�T����c�1���#X+���-�ab�#q�Z�B�{\���z�_�%�B�lv�Սa��j��!���z�E����D9~0e�rL���[m\���13��w}��@O��V�A��Gf�$�O�y�������,���������$��������,�,�?��m9�,�zh��V]"Wk��aŜ��k�k�6�e0y$�B@��ݖ�d�r��?����6��
�8���BQ���+���se�O�Ma�EI8� �7`�@��G���,f	A)ԋe^Sd�Kߚ;�r\u��|���-�	X�c�K㒙\��$uN�I�06����!��Z���f�哚Yꝫ��_��&��n��a����!+|n�o���	O^����]��Z ��e�2��q��N�0��3���ӑ�K�k��w��������V�7�U��m3��|���5��� ���:����S���o��ؽ]tO�#%?&C5EvM%i<����Y1g"#R�iIĨ�Gͭ�8��i�$�؍���n�b�HԹi]Y��� �ޓ��K��ޫ2H�y��ӄ�lA���S��1����5i6�����|�u!�2(���&��#X�!0A��!��T*����cjҍ��8n�zw¦D�()��C=��6Oz�+��v�9!��O����{B,��k��A�t֞ۛIU7}�z����������m(��l�&����Q��Շ�(aU�d¶��z�.���ἃ2�p\)'cr��BL�ؑ�g�L���3ڣ����5��~���d'"�G�gi���:z;������P�ʉ��\5�h�������d�䖢Z����r	q$r�yb69�ŪeW!kS�/H {u�{k�\V"�^dyr��	��X�r,��'����Q0e;M�V$�11����M���?C�8�L�L�s;�Μ-N�z�f�G�*���͚a�$l@����n�^-�X. ?	�蚔�ZUd'	ć��M2C6��B=gPFs�k���=W��ѿ�D�U�%��H���?��tLWbEj�T���u{@�qy�xs��T%�������BK�#=���=�\(^��hrW;Gk�]іN�h�S�?�̧>�}�>,RLF;��pS�
��A����͓���k�B�Xߧ�a ������V=�^to�l���F���ԙ�j���h����[%1T��tyd����l:4#��
�˗G�ws/Y����V�,Z��v���ܵrQ�T5�ZDfsUW����NW��� �^�Q ͺ���?�Mo1ۥyؓ�X���*(OѢ�CQ7'8�4�b3մ����7:��};�'��*x�2��n|㝰g��Yn��;R�ySb|�z҃�Vߘ�'?��]֭��5��<��H�6���b쉶�$�C�{�h�j��J�ai$'	8���
�u��4(�#2a����έ{���vq��+�#�R�,���p�����U;~s�䯞�y��K�Cv�gK!1J�&)�f��! �	�cZB��z�� �=fڪ�m(�$��`~/E]gxzV��� 	���Z�~�v�����`�*�^�TW�[�v����>�s�A��V�ܢ8��6�4��'��v��h~��g!�9����tՀq+q�;��f+�}�V2[C�&I=x&�&K�V��E��O���������� ��o��ޙ�T"Ez�J��4h����M��r��40�W��l�M��<����Ը�6ۍI+�M���O]��p*'sb��9<]��*C'�m�=�6�!��<6�|�}XL�NÇ�z���s�at��KV�{���le��� ��?�z����^��	���W[Q� (kő`����)��՝:�1ZIf!0�����b�� NiɈ
�i�1�{= �o�U7��B�?׶PQ���?s��U]����`]�� �C�^��-�_&�M2�1���(�~ :���h� �u�]����EO�4�����&�9��A6�����E��A�א��� |m�5'B�R�i�L�@�v����n��Hz	�� ByR�&��X��a�k�L�s�lA�׻���Dx*/Z�OG6�9�*�O�q-z��)����s��F��8����]�h~U/^-����e�c>�<�9̵.�FO��jF�v�uN�$Ř�XP�6gZ����,�v�ۇ矻8��qP!k̆t����o����[*�����X1�!K�D�{#�cNUc�)�,h�hvos�8	��3po>��7c������O
ﰅ��C�������-�����}}Ά�����q���]���0�EH�h~�b���K�[�������"�ᕈJ]����0�9h��苶�ʼ�bԌ5~k�h��l2�&4��]�9���̒�1��^&�[��u�*G+�m�,.�W�m���SV_G�R�ʾ�]�s1�~MB@���,���(���㢒�)9�kS6��{�ij�~]>��`��j�����5��(���|SM�5��d���+�V�p���>�'�1]��W�A�4{�`��/��2���co�c�����)�.2�������]�F\_?�	�����5���%Hհ�JP=/̨ϴ�n�M��)�B�<�v��8�uŲ(w��4�E M���)�j�w����g������n&����Fn��;C#���3\�uy��'$�rE�
��]�8�(�~���	���H�0�|�^�e#�+�E	��[�J��"�{5OV�"�]��P1e:d�����"�}�Ju��a��~M�0(�������y���0�ϼ^��,?���1��~@J�L1Q�"����x3��:���+�����J�.���?�&o�D�Č%�LǨ�	�W��Ԩ�ǲ�>6?�J`��G�$�QN��@�S���f�
��0t��T�Ԟ=q�������&�8�����e��)�P�b]�[���j���H�����c��P�Mâ�F��@��$�[��^��řڗ^�ӭ��5��f���>H�S
���2wy�˭���>�-�c-NȱA�[&±��8u��F�5��ؕ#m�'6�a�����:�^�)�Ტ�n0�{$�_�+I��c��d�-�5I�(��m��g��X�]��z :�ץkG?Ek�<R�D���t�<�G��1�2�;|YQA�&wӦC�ˁ�x����<WWs��?�>�棢��~���,ʂ,��EpW�;�C4d�H����\d)L~��5�Vr٩�~���Cl�WLK��B��h�9�,�I����R"t�Ӎ4��v<��o�b�R����5�K&����2~?�aN4��u��;��#/����ܠHǇK��33w��wDZ8��۾l�����rZ<^�J��%)�K@D=���0��Ãʖj�r�.!�s�Ҙ%����i0dcN53y0/�&)ŗ���๛�ݶpP��o���$��46����3� �6 P�d��A1v[V�<:���T���ͮ�5�J���ƥ/>c��4� ��	�W�i�4�[2�Z<=��k�)��݇x��ȥ���{�!�5=*�Eye�֬.�Y��Eb��'ϳ�6B���H;u�)�84�O;�����H
(�(��>��5o�X�]�����y[+�p qk�$MI�m�n��Ԅ��E䰴̷���$����v�,��=�h 6�|���̊�+s졦���?��AԂ׼����` ��A��Kaêo�۬��K$��
�9�LҶ=x���=n�A�$�j[9<\���O
z��gG
�M_	�Z)Y 9?~},����(|P-{=��o�(��a�ٜ�NzS}�j��[9�>AGg�[�
i�o��O8,�f���#s�����Mh<J�S���k9a K���F�Kg�w0���[r,��y	Aau����T�z(�Qc����`L�L�l[�6��{v0�|QH����f�&yH'+��|��
sM3��D��&a���qY�������㋡$��6�/t{sX_�2­j�q���	6L���:�:�j��: ��S�	�W��(�<�n� �w�?����Û�[kso���/$]��Ph�Xl=��H|Lo޿�d�g�Q0x\	2�0���$��9ez�ߧ�<^�2M�V�� nͳo� r�眈�r0$��*��Ԣ���G ����#�gSd�ҖǊl-�9��~��]�	�j�p��6�Y�Q��~�q��c��L ˙,��3�q�x�m�v�%TZ�+���;��j�8����+o��R�M�d���܆��
+뼭9c��*�~w�ݿ��,�f^U,[v�c�nx������"��?8R�8J[ �{G���~�%�P��ʐw�5��IC-��-ӝ�wU�;X���I�7ǁ�T8?�;^��(f��g�H{hL��[P�����?�	�A���r����d�Dl�����6-�?����R��n��Z����[-�E�ے�/υ:��v�d
g�|yzr*�#Q�th��� ����5U��	��	��(���?�����*���k�F�^�7�&ȶ~z��f`�\�&������~w�O-ت��������g���W�ϰ۩U���dBb�3��FCn&�����r7l�G!帟i��ŧ'�]f��:������)ёs͜˂]������2Ro����&(+/��UZ�����)9T�W�"[C��u&���<�2m߯]�֢j(��-�N>J��GE�E�-��g�>�ٗ��Hܮw��j������QxPM���{��E�86��G�L�Us=0����_	�����C���w�Ӻy��/߅\D܆�2)H���s2��8Qy�v�֧�<�dZH���:[���6�Q��U�z�f�j��iT��U���P�n�9�J�Z43������"\���>^��d�A�#�|\�*rq��qL,��c�����'��jE�W ��ư�?}�e\��cŽݹ�|@7��M=��W�q�P,� 3 =@���tF�"�<=k�y5��OXѻ��U�g��-Y_rq�a��}6)쥨r�ڽ����4kM��-ʝ �e��v�a�`��q|M�t�~�iBSAG�+���8��D�
��O����E�"���,�[�#����m�Մ#�����(�l��uc��pSß��yTr��l.ja�D��BƟ&w7�'%a��W�_`}K����*���;{���Ww����Si�8@�Ů	K۵����x�f�B�8x��3�uS��(��}����hjx yj�n���������� \������z�3R˸(�fSf���k��T/ ]��D�¸ʅ���c�>�l|�䐚%ݏDKp�տ�x��:k���I�P��4�4x��3�;n����*���/�����[ �(���`ֆ�"���ߔ�&p����r�j2/��)���ju�/a���~���B��voܽ��k�k�ymNq��5�3I�<?����GS1�1.Z>�� �h�P#��ut2�>��B�x�br�E�tI�۪�X	����=!��V��nh]
ѿ=����wE=�'yӦu"t����cN���if����
q���J���y �|I���h���[L(�~��)���G]�m��719��!7�)����*I���E�t�z[���x��$ltY*u1�`5�G4�����%$������PP3+FB��Ɛ�����sg����<��ȑS"4\>�����Y��
V�x�O�!١[���ީ�w���`�,���<%EZ���C�(�D��Jo���?[蹫��Y�ڎ�(+A4)����3|XfJw�1S������&�&��ԏSE�b4j�<�dDgz�)�
i=:�)���rf��L��jX�68��}W���^tn�)��5�����z"���a�������������g��
�dEV@��L7E-��Ru�^a}�y�hoC���g��X\A�D���wz��z�A�q4�ͶaP�0�aE���|�����ˑ���N��p�O����@7�՚V�q��Qm�/4�	3�7�^���!m�}8P:��v��."C�%(4-��o�Ւ���}�/���R���T�xs)X�`_l�y�-�ʛ�'{�ٰ�������S
�8Jܣ���Bㄩ֡�f� � ��5�G�r�7�Lu�0ʂt
�v�+iB������F4KJ��L#ּ�g�$jz��Rf���Stnu.�;�JO���M�\p���΀"Q�CD����I�8Ѹ���o�G4d!�nKy��	����t�Î���a+{�i�o�;!���n�?��7M��� J����Ӌw3���eFsX��↦(Cw�!pr���?$��1	��d���E�~��"q2�P (�˗�E�*�$�= �B�u�����Y�GNQ����Y$&��PN-�ڦ���W�eo��DI+�x�,���qV�a>I��Α@��dt�!yK���{���Z�~��pk[e���(�Y>M�J�X�E���GB;x�*�Ih[�m�$5���Nn�g���5�/�"}�;�QG7S�s�K5�0��٥���a�+��{E C�_� ��I$���<x����|B�m��g�1 s��v� C��HWz���D�r��h,iޥ=Ӏ��΀[nIX �8n���+���h���8n�~��O�5�m{��^����8	c*v�B<ɽ��9<2H��-8���7�؛���s��v�߅��*8�W���LEӿ0. �ܜpGt]�s�Fz]%x�9i~���/c,~#0�Y�鰠^�y��	Ѯ������Ҕ�
J*Gx5j���*�,"�f{��sX�%[z5�?O���D���W���k~ �k�Y�s��s��B8��%'1�}p�c7Ѥ��F,1��F ��yIne�P�V!��|a��0D$}��?nk@C��O}W�}���q��WsZ� ����TY��0�������x��������e����0Tۨ�$g��37߸����k�y�wVk��ؚ�"��9���r���ڑu����E+��2�,����>��
�z�ϋO�xPfȦ�"zf���F�o;�����>e c}:�R`�E�[lU��SN���2������N$�1�����Q`�Ծw;B
�/��"�i�
�nt�>�h��m��"u�e���W0k4�ۊ�VNv��o!lc3�`���ޟ�q�U���#�5�:������w��<�x�D�h����3/"z>©�<��R�3�>w,Y>�6��P�*U<v�bW��^�׊ʈ�!4����Q�����(L�wS��H��L9�	�P:�4�hp�z�lL$�ل+��l�"׵\X0�R�~��=�P�I�[��.�
�<���9p�q�����j{�j�'y}�[�֟[�eN�7��嵚���������k�H"}�4���SH��|N`
��\FC�L��a�^:�k�4���� ����.6�C�'y	=-N�r^
zN=Y8H:p�ċ��3�O��x�ڨ�ͳ�H�kAYæW��cw�Z��������q��].�5_�1@t���%��qp-�a��Ig5�l����F����� ����ޛDoI��P3\\�M�^��"����TM�σ��r�2�먾v ��^IO_�ic�~�R)����6&0~+"���q��1��Gu��]��.?��C���ӐG�ۏ�%�e�eo�����ا�5���ˈDzL�����ˈ�	����p�J��.p,S�EG�N��(����  +	\�j�}7$���n��ĭ ��)��H�Ʒ�.�ui��7p4#P@�)!��Ү4X�Z���".��*Ԩ�
����Bf�?�D�@�ז�z�xx�����u�>7 f7�4:H,;�m��ݶ$�ڧ�h$=Wi�/�SA��mS��kq�����?��~���6�_�����'��	�}R�[ob˩�W�g���_c;g��?bR�z��8Ʉ��Ak��|c��{���L	��2�c�����!W�� ��v� <G�6��,Vmw�;w�8m���6�y^�I���I����,$�d������I�bPO�&�"c2I�C��g�W�A���T�E��Z�����&I����l*�X٦�t̨[�߭�{Y��2ʹۜ���(xE�iݧՕ�w^e�j���I��ݙ#>d��SD�Na����w��C,Dw��X�v�C@W�/^~�}��#5���=�'��#J˓��UЌ�7M����z�V.��-q��4R	��)3\ X-D����~�]����3��U����?�۳�R�UXD6��NK,��[:�|�T3��|>�fO�x���M+2A7h��Gcݱ�Nu$.t�\G��������0S�ِ�s�����Is���Q��:䣭��U��9�F��+ϭi[g�J���a����0��5j,�|�ӄ��52A�P�|lא�BIbo �)� �=��\2�5|m�f�j��V9���>�����;>���
�8./̓�#]@+�M���A��Z34�!���v��w��ؼ�c��=l"k^���(��~i%��Q�?�学O��W���\J�$���)��6�+�e0���#� ��]/����l�����v�� ����	J �55 ��mM���<�Q��I�.�]O,��� ���D�8#�8��%�t�o!��'��݇�|�!���x��r{W����P���Z�����h�+YXf3��=#$hu"��ֽ�0�
�~x�)��!U�~�T��H��%�/��G�C��`6ۥ��I�d��ǌ�P�\H��O��K&��
�h��)�
�eZ�؎h��|i6?P��bS��`�,M�~�;�5��ԭ<��P�%��8V��i�1V%{z\� ��>Ap�=�܈�F�>a�0Ǒ���[jC�����v���.0��i4��Ix3R�j�=��=�ıѱ�a ��L)}�p�jDX/=�NBϕ6���Y�]�I�����Fi9���_�)Z����H7��RV��������|GR(������Y�$/�}�xi�
�G�<r�ڨmh'0b����5<m�pv�5}6��J�d�ZZ�.ž���m��� ��K�q@�R8aUʎ�>�JBRb�_g�`�,�pJ!(ӭէ�'yW5;����*�w<ݏ}������"��KP�Џ#��M�Ŭl�M��_�o�Ǐ%��a�eAl����뇿/-�*1�ui�鯖�_o������	#�KvC��$�:��wG���CI~���jz�G���CJh�%�w�{#b`�� ��E+KW�~K.6���c?o��ҵ�ZyY\�;f�I��NY�ߧZ����{�!�h�.�v��lPYڗ:�J�؂�w�sC�_%�ߨF>,"��������D\gc���"�'|~#@B6y��J�wS���`�^�:�x��z��ma�������[[� �y8��,�C�c-Sf�V�{)ID5��U_l:�猛g��|�����?gn�LH��
���C�d"�6�o;gHs�8�TmU#��<r���>�xۺ�>0��LL�����M�gd:�~����)���h,d�womԁG��V�w޽�T��_�ŏ(��/x�5�]�Ψ�D�����>lU��X�aL�w>N�xՂ|a���z�l����b� @�y�`�C��G��,�a|摩8�
�^�����Y�'�b9t:���)�F5�=�C��d��\Ú/P�.�����/-�P�wш��,?5hl��~�-�Ǳ�Ma�!v&���ی�>�-����$ �����=�����E�n��B�S�.�E��݊m�1�Ğ�x�<^C���q��I[������z�:ɊGW�Է���W[�D����I�^Wl�k��N���+��W��y�+�D!oH���h|z��p�<�(/Γ�P�c�dQSg�L�}l�$��+�i�0:H%ce��j��H)�UU:Nlq�C���K��p-U�l.Į�1Ur1�T;ze��M�*���p��2V<�5�ڃ�r�>�A�K�f@�U}d�޻%Yˡ$��}j�B�Y�Ԝ1
�j?�8Үj����'�!w�.������J�	�~OCٹ�����jl>��O5�eL"�f�:� C&jf��#�)5�,� �vu�$K#���9�����	��b�=�3�AI��Zm�s�^�T�1 �[Y��n��1��b��?��2��� �����㭋V^����q��p�No�T�M�����ACr�]��#�*���3sJ�o�͒�	��t�۵W��	Q� �#iB*(-,HL\�Tp��|x���߭>x�]�����A8�L�Gi�k�j_6������gIH$.�s���	W�<ZSߴ���i�s$GhD���@���?G�^-��a��M��\�c�kZ���9���V��Y�������'�n��i��k&��3ӥZK
�(��\v��f�{)�f�`�U��5���
�K��c��%(�\���1Q���露�P�Q���&;�x���,��=}����m�k����	� B�5\�!=��������Q��ޙ�D�5~�������̀y�!:��<޵c&Gw0�{� 6�MJ���3Nf�L��w+t�����P�>GXi����Pm�*m9Qy�TW"��m���a*�{�NE��k�3��)������ߏ���k�����u�����`m�fMK���b�]5&����]Ծ�7%������=����0��`�&TF'�@���"#õVD��riR�����CtVs� Y�i2�-���z�O��X���}y��(�*T���%�ʛ�"����l!�v����(:�IKߔ<h���vYX��,ܒ����"�;�χ<��aWDx�A��9��ѴS��f���,����b�ύ�� ���j�?��m�e8��E&��v�����:y��:�.��o|���GC}�D���Ҿ\��m^S�{�� �ݾ���>���{�gF{��'/؉��!˹J���ȑ[�S�`	n�C<_�O�	���ȪKG���B��k�D<���� ᑣF���V��+h�ru�4U�[�47���������;zM�on"���/6��������5���˥���ƄgH[;K�~1�e��o��9�o3� {��a�a��G�����.��sWИ4ϧ���[�����q��D�ڵ^�
�p8!���\�P(�kңd`�:O�9bE)P���H o�R�"�A�9-�L�`M��;�(p�}���l �ъ�:5@GǕ}�_����
��k4��G�V{����/�S�(yZ	�=�����9���˹#a@-;`U7���=DW�n�:.�K�#�!�|/YG��.9��_����r���ʛ����F~�*��PrAI:�̃N�����G$~����_��
�w<-�bl��~u�]��ɘԿ�.�]�E�s�΍�<i�c|؂��(���m����Q�J��U._^�L�&2����(.�����!>R�m���	R�p�Ŏ�����a�g��'#:�еK��\lN0�RI��x�eY�������B�T>�J�/���c�#_��t�:���?t��+�*����(�q<�l�K�mEu=�M		%@���7�ݭ$�X�J�˽4&S��y\n�K=:�s�*���M�z��Y�-�����-(��'ϥ+��Oe~-:��>�W��Qu�ִ��g5�34y�GZSD��4��1>�M<��K�, ���cM��R]���"�W�q7*��'W�[u7�Ҟ�n(��w�h�jK���e���	��[\�^��`��,��74N��8����Ŝϔi�%�*��F OT2���"o ��[KD�oj
�O�>� �vN����q��1��j�w�Bjѡ��=|C��0Yt�>�q��#�H^؛�Pv'ǳ��y�̋���A�*C9R�*�׎^���Jq��]�P�t���N�*�	�)F5�#ʫ* HM�O�}�J��\�N�G;ac��bh��Q��Z���9�]4��`x�%���������+�2>X�,6����8����c�AB!�[�����sVEϖ\�K���㎆Ȑ0z��G.(��?���n.O��/ʻŝ�%ǎ �T�L�-v���QX1��G�Er�o�y'��͠�Շdh��j,��49k��"͠&o�F�!�͛�41�k,Y�df9+y�o�"�ŶF�=7S���I�U����c+��ՠ��_�O����&�1t��w�c���2�m���ҥ��o�'�ߠe��"R[�����b�k!,Kfц� �"�}�x�,<�G�s�K�J��%�aooQ-�t�f����f^�� C�b�$;T�3&)���|�}�]F�iRp��[�J�v<��)�NWA��H1�i�
'F^�/GuD�n�L�f�v`�ƥ#E]�;CMlYh4W��s��W����sD=jZdóx�8	T�*�"��=�5"_������<ˋ
��y��K(�Lɨ0�T"��T;����j��n�11��A@�����26���78r�>k��c��ay����YS��.qUl�Dg7a+]onX�񼙡��Ւ��=|��rZ6����,��/���1B�&2���@�g[��MТ2��4�����k���բ,��R�9D�zesF�u�nr��۠��Z���O�����Ջ*�éB� 'w�o�~�ų6��S�X���T�����1��;�+��^j�6C�Qz���� ��搘7�mq����f���C��b.Ԭ�7�l���q��]B��!U��_�3<9�s���7�3"nY�+�_�":�gdjNR���,�d]�L� *���za�x9�ҁ�x��'���:�na;؃X�V"�9@��Ǒ�B��?�{���u����	'5�?\�lK��[�֩��g��5�e�>������M�S3��={�ȪyrPйE�QO���Ռ������9,�E=���Gɳo�,q�hDr^�F��aL�;s#@���{�������o�����m|�S�'�z�H)��A�Ԏ���X��Q0YMP|�~^�T����X�^uل��j��mb5���*�������ЗiW;����������X�˻u�����RG�.<�;_:��I��\f��e�L�J	�^!C�a�Z�!h<�#�&�K@���7]w[��������g�Th�[�����x>��+�댎{�D�q��!�	`�Y�w��n��LD��};���Vd����7dL�όH0`�����E�}�ԙ�7]���F@E�u���[��J�����Q�<>�$k����ޅ'�!1�)q�����b^1=��@,�<�Ei�ݶ����)�Z�=�x��7�b�S��N���͟�g�άʧa+���@ۀ[z�.�W�Ŵ�i�#k�9z��]�:}{��'9gX0�����!�a�=�Ș�z��
	�?a?�6���/��L�}{�փJ����&�p\C �?@��%2��Ζ��o �sɕ��)�w~����:Y�����#Pٸ���,���?v�dy�}��u"�xܼ����Yd�Dm�Tw{=�e��y
Ywop.��9 t�H�!�w�qD��G�/_�΋SV���#�H����:Ig�!���3O#���=OKU���aG�㲛٪�B7�i��V����FS��nktL?-�����L����֩�k�mUQ�Ν(����1ќ��1���-�*�:��,)�E��B��`��Z�I%=�$\4�BU��L�/��n��4��G6z�x�(������P�s�c�|�f]&���>�н�E`�6멵lsΨ/���r�O����~���ձ !^�L���E+�D�o6��4�s�
�Xc!����ӣB,�� j�f0�����W�u�����cd�8�c@�sF��S���,������D���y�^�sC|\���[ԫ$T�͑[��ŔD�,�Cvϙ�ѩ+�Ϩ�����]��5���(�[o�qIq=ߟ�i�:
\+g9�Me��[F��H��U��ZDc��tq>\W����I�0��5��B��phuXh�MF�s�6�yɋ3��x���M�k{�¬�zD������ﳗ�ۜ#�᳑�Ĉ67�Ň�&��-4��2�&��� Gq�s@B[(��q@
� �(f�?��;1�i�G���Ƭ�=�����2�*XQ�']sE�w�����}؂��M�e!??-��6!^0"|,���>K�]g��&;|�l�«�g�,v�8��!p����3��ǆ�\�wx�P�>�]"4,��{��q�Gɂ�<�s��yR������������b(V��c�š?��x���~��\��U}n�k2�\u6NJ���}/h�K��z�i}>0��B�Nc<D�֚}s�'����q o���*8�����r���ʴH[�[SHұ�X�1|�����VI�@}q_.�j�1�d>��m���T�ŋ&���bk�!�h${��o��..�~�V�D�.����4�N)b�����>n��||���kS��R�Q�fDW��
�c�q� ��I��JI0��_�W��_�v��F�`婓���uTQI .�
��i)��K�O�%��Lv4��� w�����t^W��
,�?�N(��nSa�+5�B8$Ǐ��G���[sVp��j�{���1:Zu�$(�L�E"fU�;a��V!��qǏ���X�t������ C4�O_�U�ٓ&}�0���ei!�y��Y[0^���Y����8��d��v	����zRZ��E�E���T�CC�m0E��"-;�o�e|�-ѳ�d�L��<��ݑs81�3,F$��H�������bOy�`x�c[ΰ���}-���/&mKq��7W棕��Ȫ��]n��K�w� &:���rd�{�p��� o�LG���X�S!���J�]ٰ0<U-�����9�L���,�R[ߋ��`��p�N&6>�mBm���  ���Vn���-�e��ؿ���_MF��A2��l��gR�WͨB��q�#�8Ր6	JU72�(�	��������5`�r��Q�v}`P��b���������ވ2��-��l_�cV#8"�v�"�-gb�J��#ߌ��O4ɑ�]'S7��,V�?���s�8��;.4�����ß�>b�M!2c�3�!��{B�ђ�S*�HD����j�7�ؠ����"gj���K�\*�t0����k��\�A�9�v��+C4ha�s�#.�����
��c��3ڨ����ݴ��H˔G�=y%�[��@[G������B���dD�#)���v�R�����_z�nz��N|m�'����V�Až�GjٲnY�!S�IyeL@HA�9��w�Y �A�����lD-�x4�:k���?�/���X?)�e�r�n��UYw�o����|��;�݋o���K�w�b���Ƥ��:ɓgDy4#�f/�����2�:��o��2	 ���i)� �q(�Pl�x�����,|��it�X��x�o}CYƨ�6�Y��(������xO)��YP��.:�.� �$�m��uz�V�*<7�F?���5�3�9�DgCd1�$�o��@�i�c�&�:����Kp�Sw��a0T��O���v~�@'|ZL�+G$֪��0UЧEa��)��� g�
��:�w�; �)ٶ�>�8�V�R���Y�/u���_O���nښ%9��P�e|���	��q�?�DrGY%iX)8$�+�� ���T�������/QY8��E]^�
2��;�����,��̇��d��#�&��Ix�ψ����<g����.!2qW��'�_	��V�OI�y�{)֣�����9���ʎ����Ü-~�w6�H��I���hDEn�g�����5J9?&�4J�s.�e��kmiQ�	W�8��+�J��E��1ܴ>�g�>�eRk��##�)��>�
{�M@`T<�K�8х�������l�l���ٙ�\uA�-�	N0�!�岋���op	s�NU�7���J�P�q���Ǎ�rMt��l�.���Y����)���������W��N������f�� sќ8���.���<w�_�{���0�!Q
�pm����%���{���NO�^C��i�S��HܰE�w|r�&�+JS<�Μ��=���.�K��3PWQi8s���~pn��޻�P��#�iS���u�H��P>k%o����`��|���,] ���Wb�O��Q���K��W�w�}^��Ѥ����J���!c��qL����������>��S�\����R��r.��0e�X�K*�!��%#p|�lf�-=�O)��l��vcX.ST��5XldV.e� h:�}��֐11C�����Ć�M�ד2}�b~�Y�`��9�����~]������%��a�G��m�ǜ�_���
G
K�U��7��.8����i��:�g�qr����	���6���\r(�x��w��i�Ih+�(��1���Ƥ��,��`��Fle�U�x�ur��	Ɖs}>�Y���5��,���!���o���4�qE�%�ކ�-6J4V���S$S��6��c*�>��)�o/n�YC� ^撽��J6�x&�^lI0D���ـVX��h:�A�� w��\�p�2ß˟1#�r��(��
��La����`~�J�l��E˘��.�HC��7��O>�F1[�+��ģ�a�Da)��LT�y42)>�=�ApQǶ�}��1{�l�ƍ��� t�?�{F4���y�-"���.���Cj�#jh����Y����A��U��5�(d�=�<X򤘎$�9�i�F�m ����XI�� `�����щ�	�x�#�N�A@r��)r��ªO�wWiahP\�"~qnl'�eJ��8�z��G^� ���(�;�TX��q~Zִ�� e��z��ŉ,���O�gV��حQ���v���^��bw�x�>�kAt����sT4��� $_	|���¨���w衆���z��DyI��T�� g�֗����7,�V��������|�c.�	;��C�fI��������rЫ[�.�H˃��[T�; ���.ˡ�C�����r1(�O9�Ȳ���-���0��L�+K��Vm*w//-�13XHM�)�o��"l������2�P����y7L�@��lҟ~�o*�~� ��0R��oֵD�N> ���:��Y�c+�X�P^�x�z�����-�*���}t���ܢ���%(v���-����5�����H��XԔ�z��]�\E"�X����i;��]��!�#})1�#�e��JI��7*5\0�O�V���^ݪ}��L2=�	,��8ל�(�loQz��4Ş��U$������XD�3O�D�Z85t��y=�J|��7�X��.c{����rs�L���5�%���K�nh���9�-��ZvWb(FU4R�@��̀������H�r�I7%̻,�e�$�C+}+�d���Ņ�L�b���ˠ�]��7:�Z����h�,qR1�?�|��(ïl��yq�a��j�䩎��t�������Qø��H��k�^�BdT�$֟��f~�o�.�V�(v16�54f������fh!t K������a#��R<*{bh9����󕅖l�x��-��/&;J�3<v�-��%`���o�}���P��Ѹ�ۧ��-w��gr��z���"��p&%v;^�&Ⳋ��7:p��W2?����qi�K	j�c��L�]�p���R}|�<�q��M��E�Q��3�'g���IV}�^�S��\� �Ї�kE��VL�Ndţ�{DѳU�8b�9ɞ�t�Nl��*O�$�A�5�Óq���k<���m��R�F�U��mea{"�ѣ��0�gn����	Q����5L���s����U���߄9h���b��_Fm����R�S��C'd�k�����Q�$�*<��g,@3E���K���K�����Y���pq�yN@$I���~ul��Xvm`t�
ٛ{�V*�ix������g�a:��Kjo��i�o���Ŗ��C��3���8�����Jo̔p��[_YuG07�$���)��:���w��nG��+o���_���x�E\�?�t9xLG	[��N�5 �hs��(eF�9s�j�uy'�g�G���Z{��FCEy�����9���ZՐ�w�Vט%Q�����)����U>��|Oe�*��m�!�ll��_��Q 2�y��3KAS��c~��_�y�Y�����մA�������	��{�t���M�Pl�K_�Y�Z��4��f�f��������������+Q�T�O��h�ۦu�f�Vqi�|��������g�f���0���R\IlP�&��>iE�C�=$vˢk2?$"2[?� �k�ܑ�9\�:{A43����cu��7(����ϖ蝄����\��qZKs<����8��p~7t,��9�}(��Zw�K<�p�� �k�{�4��Jvԥ���|�~y�`wɂ��� �~��)D�*݌�|�v��[<5Ĕ��j0%���X�5��˂���#�7�.:I��H��pF��˞,����o� �gF�K�[��	8�.������1��Q�ϊI��ހ��"��Uu5��(z�ؿYr� F��bJҚ`�k���\�0�y)/w�3?�R�)�e)j���=�;�a��9^lj��U��<q�G�|�� g ŉ�u�^(t�.̓�Ǧ߆��{�����R�
�K��;K���S�ʝ�?hb���0AO O�u"F��G��M7�ˈu5�$�D�&��h��SG���0�՞P4Ia.����o7������^�@�A�I_Ly�n�H�����y+&�n(Ԙ���B���k��E��_�<����c7C}�
���^1!P��D��K�Lp"�z�ޜދD��v�F6	�L��s�wu=������e�g�.�G:�9�Й���d�1Hu���/����@Jň	�l�����g( V8��ª٫u !��{��eY����?�O�C	GG��"0�E����q�ܵ�Ժ�G���"k��,OP�u��=��ܴ�׵W
�͒ױ�kx�d���2c.+7P�|�{�\>�Ш�O�w�,�N���ӆ��IKnHW+q
N�SѳX�u{ޏ[�������-�_�!��5+`���M��D8Ȉ�)���J�����_4������?�������NO �%�͖�_��ٍ\#zT��@P�s	/`��&n�<��3@�����Ϊ�m�Q�E��AHc�b�!�m�,`��.¤֝�x6X�g�>ɺ�OZ�Xv��)֘p��:�+���)WXk)�l�Ġ%��$w������1Y��DTH�̍�F�P����nc�ݲ�S���ԡ(e0<���a,n�8�s�?�٤��_G8��2�*���#�t��!WLݾe���Ř�2ϛ��I�0/s/0X�3�U`kF�����^2�s��Ň��)�����F�1X'j�!���l�1�,"���z�B��`���VRr,|d	<�h��ꈺ�jj�p�L�_Q��b�G�t��T4g���?��Y��D*�J�El�1Hӟ3F�^#� �'�i
�+r��PdyU�_�H�Y��%��s�OG�ħ.�y�)
_'q�5���7���m;o� c��T�W:�U)���\�J��p�fE@�V@�x=u��p�c�2�*�`��9�_�s�
��V۴�-�k�����Bb��G� cŐ����Z3��J���A��=�����I��Һpb�qD�W~bY����ӊ26JX�b��ҥ������ı�וg[[�ꭕ�x�-眫[~���`X�P^5�}5?�p�[oV$�79����{�&�6s���*��I�z�U8��l��Mb68̘��� ��.%�1g�v��X9O�����#y�%��\x�B�=W�A_o�ZxF#N%Ϩ5=����Dȸ��ȤK���yZ��m�o<�w޾d8�A�	&�i�M�E�u�i@OP<�Np^��D��t����g�x(Ff���o�X���i�\�����nC�Ǳ�c�f.���/3E1�u��ߚM�d��s���w`���PAZ�v�����|�TO���:S�_Gl���hB�\$ө�ٶ�Tc��O�;l�L�d#�	>��[g��´��J:2yl���Q���}��a/��Z�������3*�Y�W6�K@t32��ܬ�cS&Tt$ծ�
7���ϔg�ٕ�v���*Z�|]^����b���dp�}�����D�	�W�Hs<�iJT��.W�џBap����Fi�l��&nj�����	���6�tP������ D��
�9�J�?�9zN�)�Zq
����p��0�%�^%�s��fkY�p��V8r��)%Yc�YE9�L%ڋ�{X�I� c���d�Z�u8� ����qW��h�b�1�Tת��z�ph�ai�9�o����R!��d����W�d��?����r�\Z�TܴmñH=����iH	��,dlAo��HM���2�AV��c�nX��Ž�����+�~�w0�k����H��x�L�'�����^��3U�������f/�Rj@�;�^���;HR/�oG���׷�]��� ��]�p�_�C���w \˫nmL���!�|[���(īk)h��ܿ(��qE���R�^R���Ig�w�w���P��W�c�����hk��8��Hĸ�5�S� 7KaX?�ϕ�sN��B��	��o5$�w%�p�j���hY*�X��� Bi�y��R�jC���a_��ε����zĄP��y���X���b���:_&)p�N�5�4���x���EA�[/H�"yg�=�^�$C��55��j��m�}ݟ����pm���R_���R٪7~b��I#�
�y�l�#�֣��������V�F/8qpP'��X�0���cR�aQ�l*�@��^6�%�ށu�F��K���}ﱢ�|�&<�h&�E=O9�>���n�*��/��f���Hk�q�@�L`0�"#<�/�َ�����b����o����,�׾2�7�H�8+J����G�u�_�x[r��(��'!R� ��1D�V��g��h�۲/%��M��`���g�y��9�`�\�x#�d˒�����tPH7��?�y�ÔD���P��2Ңoj��'�����:M�eg�_J.)^��b�_m�?-�'J��G|`!��ŭ<���7ߗ�����F4ˁj�,9o�0j��I'�7mH�H��ߩA�/%5�F��6>|�C4�D���]��I�W9S%f

�6��'��T�[��2YtK��^g��]�:�¤�V���k���_c��0��!��*�2oևg-/�40�-���`���A�� �c��Ւ2x���dO�
��O|�<�4��[�b?Ux:dEqTD4,����U��/���r�ݝ"��a������X?���O1*^�	�&�1I�RZG5�茡��T���� e�L&K-c���x�sq�#�sө���wzzc#����k���*7��֯�m=�w�"��#�+�Ge����6o��IU�sC�.h��܀Y��;�%|�g���9��y��c1;�Y\�4n�LV�8@�<ȝ�9��<#����Kǥ2V�G/�?������
��E�J�0ݖ
Uv����<H�/}Q f��#/�5�Vĥ_=e+u�v��6���)T�TR�i��̗�bW>�pQH��k��h?�B�5r]�,܈���I������mk} Kؽ�E[�\h;)~3�^iB�s���9Մ
�&��L�<������%����;�{^x�$��I�A�D� #�x�ԋ�WJ�7>P��N���C3��0�1"*B4��X�ޯ�d71|�I����7��k��Ѐs�H��S�=gH�5!��y�\4��_��; ]���|�� K�Y7~9k²Lu������)���Z��� y%�53�:^�W\�,A���1� �<�>q�9=z�*-- ��w<Q[O�;��>XKg5�點F��^�n��@A�\k���M��J��Dge��07�B�
��t?�7j���C�%� ���zJd��d�]�cB¢GO\���s�E7hJ���'K��3����z�(�4�O	�M'�50刕D�eUJi���T���}k��Ȥd%vEr���*�M\��X�����
��h����!n��D�c1/e�.�����8wL�E�3|�ժ}���1��E�m+A;�zs�H����������§�Up���XW��E����^({I��7��d�Za���>w[z� ��T��nφ��b]L<U럕�N�D�\��P�<�G�&3�hŅbc樓/�i�9m#�S��1a��9�*V�:[:��#��Jt��f�w0C��t~V��6:kU��2oiT��A���L(I�	Z����S�lґz~�W��ϥXv{?@K�t��u>geP���/2������Ǹ����?���~���L����+w�q��*l�s���l�urZ|��
�zS��}��T��R'~���й��{�� N��������C]�#]���cqx8;��=N��m+�Qs����Z�4�%y^�!�f����[Rn�G���׬�e�����w5��0��SH�e_�~��2���b<�w���:��y��U�"
������,�����'���t��u����{�2���8��
��w�����Oȇhk��-�W�'�G��DL�:ET���:R�hn�!��_���%(�@]��1�	Uˮ���5����Y��L����4��;�ǳ�sAMT�J3�A�ԯN�y��G���ZܙӸ!}#�E�r��ٵ�ˉ!Nd���.��&=193�G�7�9�3?ҧ���	k�Ęw+�4�P���8��QU�ݩC���n�f6Kl�on�:!�n`jF�|�ws�_x�u������iSL��Ӫ��xCZ�-j�����Q���� �����c����գw��B�^c��h��49s���{�5tp՞{5���Gq���oMe�LwoB��X��C���������t
���9�C�y �~��j!���c]JEYo�*�_����?]�6�w����=_�Ɍ�1#�#gCc�xo`���up�j�A�r4`ETϥL,�2�#�4*���|=뽜).���e{M#�+F��.���(���=߮�tjZ����egz���g�s��[2G)�7d�e�d�[)�a��9�0T���* �t���
��-۞�[���v���ʫ�?�2���r k���l�,?��|E��I�����5�j���zZ!��O�#��jAq��Z4�o��/�<oU���v
�B1��Go{���	Ȩ��c�=bp{�����������ا	R�2��;ܺ��I�^NL5�����h*�!��w�T {��{��ط�AĆ0���)��_8 �f*�k}V@�c4pyH���>n&�{2�\%(�$�Љ�Z��FU�K�Wf��\^����l���;�6�G �a���.3���³+��JvF�9�xfJ�D�${ͬ���ci��0���C�P%�[oh@4/���>�[w}F^x�a3�k3��7��c�f�_�S�j�:��5��E�*z��C�H%��
[ʅq+@´�����ԢE��)aeе��6�Y�U�U<sX~=&`���͂�Pj�Y�FpOW���cqLg]�������B5�Z���)_�R!K��4��?Pl�Ez�*�CK��j�xLh�e����<���m�����rT�Ko/��8�T#_J������']#A�m�u8I�nњ�LB%G4�|0I+������b��4�:,G�����	-K�����F���-T�4[���!��WwEzRaʶ��9��h����|���6�v��u��82��E�#ڢ�L�<��p����մp�}�gB��c�-I~�F��LV��\���%������8}k���[��DDݩ]v�5Y+d^>�t!�J=�dF�abM(Ē��Y=�I�i�=�U?8s2�꧸�{�s��Ȳ��5�A��$���� �SN���|�e��J�� �Ih��@�fO�cX���d�]"˄���1_�#oJ�X�%`���h#��6%:k��1յE_����НX9U��M���>�q̔7���k*��BW	 ��Y��Q$1TJ�H��׊r+_�Z�$2!��ĽU�,��/�������3}x ,�Tx�"��4�`�-Z��Z�s�����(�&�Z�=f�$s� $�}�$T�g�Vx���~�i�b���E:�ZnpAG����\{��P�{W��9�v�/����%����5�`*1�A��g���sE��=4��#Z��K7���z=�oa�WW��#�7�Z?���w8��:�y@�	��w�GU�iy�����J�,���l���j�b�r�^��lT�����0�[�cLw&�lG��l#xD��#�a�1���7�T���xy�R�~�d%�/�����?�ݥ���]����e8L������mC���u�m�f#�cKAԉO �Ԇ��󃇶�����L�M�O�DY��	�g96���c�<�D:���l#z��]��i¨ ȴ�K��y��'�{���"=wقnG���0r�"��o�JfPZ���Y��ͦ���xj�;Q&���S��Yٻ�R��>������x�Pѐ�d�T��4u�k�� '�[��N�_+0���zP)�߰NK��Om6�~t&}�?[��arE��h�QJq��a�7�;���`\f��SU�W���8<�6�L( ǐ�F��2�R�=Ib��q�4v��R��ԃCI�����t>�P�x�&�?Ê �@&�p�7�yɰ)[����6�J���n7���Z���vR���w5�I����R�-�Uo���ZÏXC�ec��(�]���'C�ӟl6��)t}�z�7�Pm�B�.D1����ݙs��"ǧ�5����3�) !�q��zح�(
��2�J��ny⥅�/l�a�mIЋ֍&�PX���Z��`)ԣn����ݟ�&�G8>�El����9_���/w����tv�Q{b����2� w�|�n\���%l������r^�I	�xۇl�cU�T�m�e��$���O�SQ.�X�[1O�K��.*�`0|8U��$Yw� ��^��j�ٱn���=C%;���6Qa�>`�@0Y�����(�UV%��`2�w���s�J��Z�qOđ,3�Mu��	`�
~q���O�VL\,���C����Ǧ����
�ex)�s�M&Q˴�F5�<q�t46@,JaҥCpc^�I�����y�-q���6�يC1�Y�a�%�[;����p7�V�9�m�z��Ӕ�<������sM�]�E��e��Rq�cY�����}�P�Xhɲ��m��nv`)=�]O�r���X32aQa~v�u*�����*�dR�h]��-AF������4�z�I"�y�:��6�N�ĭ_���#"-� l��1m���7��e[0Wa��R��D�&��+e?�u�}����o�<�����叙3|�Lɮ�θ)֜�?�?���3�l���6"��%�! ��7��(G����<GCeD�#X�`���wF�N�� տ�!�4���K���"2a�C�P{���<���6�V�V'�G�.�}���A�;��t�C0�)�-�ղG��r^֊X���hIY�QiP�C<E]U&�Td�,.)�i�#G��*J]ٱ�_����^خx����lu
<-��Ca��y���MϚ1�mԷ2�'�>]Ws<�y�|��=�ϡLö�����
��IL��{��j\�s$Y��R�G[q|�~�ܚ:��Ѿ�u&Gg%r1<��}9|p���|�������l	(aQ���a����ݴ�E�a�j�+ʫ����J�����.�;�wӍ6y/
��7��F�9,P�T��R�u|��0L�G �a��`��'V�^���id� ��c�'���M��q�_yEt�e6;4Qա@�=ԥ��;]-�����O㌁fE�;nN�$p:H�+����Kf��B������6ǯVq^
���W����Q4�
{֋5~�w�����!7V[��9���V��T��(��U'-�?P��h]��*���@D��߇ӿCB3MV�N�K�N���Pȕ��C�P�2�	(�1�C�g�2��C�:@�P��(��4.��m��`����#������]��X�������k�x�����4�
��Ut-:�4���F	����bA�逛F^�YK���Y��`%�9�"O)�f�,�4�)?+��@Kgܻ�mW���NA��(+s}�D��ְ�!�/QE�h�T�÷y�}�,��̎u3/|����21
]�]_����F�I� *jX�L4 ��pHMښ�Fĕ�4�k��d�e7K2� '�K,�)\	w .Ƒ�{��}���5B��݂������WPz��|�ƽ�|T��ېR�Եϴ��~�����P*hn�v
�Fa���>�&�ڐ@|�N�D�#�Q��p�{��ڛ�<�z����0 ���� ���v�%į͍ؑ�p�暧��J�����ڵ��[�\�� &�v���*��5���Y9J7 �bH�jG��#]Ӑ���l
���/�x�.9�ix�LHQLL2I��}:vN^��	֬������/`+-����+L��3�����!�O��z>����{�U_�[aj\�C�aI���Ӳۇ�<����C_>�ƿx&b���d�8�Нcld~U�I�a�?v����/��+��\'~d]��BY5x�Z�m���p|�|y��`R����N�ّ���G}K@.�_��d�d5�I�!�Ȓ%��;%�;M]A�r��D�2Ux�y!1Uw.e���ֶ��K�=#W*����`A������2D<BͰs��;�# ����k-r6By&ZsL��H�g9,�4W^o���#��Z���қ�Iuؠ�0Q��F��D鬪3%J�I�qQҤ[g��G~���L��b���Tw+�f�Vܨ+#*�bB9���&�{`6�̿�������HҠ|��U���:����S�I�Ӛ�M e�*��x83};��%D�L�`sNS5�.�#�P�3������Lf%�R{�y�"���L\_,�u�I#�5��Am�b��<����t����h;bC����<�9~h1��".�NYʈ�:�W�`G��MY����ΊUu�v���}���o�"�>��G4kX�,�+��׸�k|2�dv��L��ϵY����k�}��:�U�r��?<��I�_�f�X���27*���Ll�р�o��R
N�e3��s+��h�b��j���x����s�kUkK���'���䜺d�P3Ykoy��%��d���=�M�s��EE�++Z��%BI�u��y��R��L��5+K%Y��oJHp��ٓ���&��h�T�-]Eg�{��"����TQ:��d�e�����iQ`í@�q)G`w���b6��%�� ��m�^�u��� ,%��R���m�G��t���0D�S��g��'��%y�#1��_:~��^�w:���=Ȕ�����q�T�|��N�Xt���&�����T΁Lx�	��6��J����M���#:�~O:Mζ�������#�������)�5�)`�$gM��vV*���!�HCQH�h��~��k��~�#�	#��}p;)�}dz��}�}�C��x���'ۡ��	�Wa{�$7��G-!����b��J��䍼?��a���k�0^�Pz_�K��bk����4�y�x���_d�j��:m�����[|��V�e��9�U+,�㇫�J��m���F���j��(�����t���>����_ə�ݲ)�x ���kXN�8*b���n��M%�8}�������$P	j$l��B�=�i�%�����}�����!�@L'�j��������Y��p�8�nb�6�������E��	��P2kQ�������ZB�ϐS��Xv�I�dF��E�Kϒ9�S�M����d������c�8����^B�E��=t�eb>`5Buِ�T$������:�e�mmv�I��L��y��vv�	�ny�
��w��"	�0���en�ib{.nt��Εj�>�I~�e�9��� [ ��_eP
����t�m�׹���w��P�T����r!��餙t\(��4\�ǆ!LF4���Y	��2��Q��Y��h���,9��%`=��3ǏU��
6C��Kt�?������KF�|���w6�Y�l���UϺ��NBS/�;83"���nĆ��I@m�2FܖV󓴾} Z���K�Q�b-��a��2�iz�Az�Kv ��j镢[\��A +L��}�00T���њ+�r4K/,VV_[�d�ps��>7E%�EY�5yx��2��~#le��+I��u=X���Dwcd�b,�E� ʉwu�Z�-���a�QtX0�%9�=gB��**��Wb�)/�2�\t��&��^�����Q�"भ�G�`A6m�����$f�����86Dq()���N_V�f����&���RQ�����r�_��Ƹ��+u�		��7��s� �甙�q���QB�<^�^����v9e/,�-���-׺KO`�&�!�~Ø7���պ����o�b�a���=莧IF.(_�ˋ�_"O�����6����K6�d��?��鍠���f�릮�*�%�������Xxh�O���
a_��
�ESnRa0�P;�'t	s���F�!<ӕ�t^�*���´߯����)�QA$ɰr��]��[G��9 ���̺�n���íҸ{�۱�����Lv�[ͯx~� ��1%Nj>��;$l���j>/<�ʚX�ph�-"�ɼ*$�L�B'��!�p��.RG��@��E�P��ޚaj���D�x�1��^a�*��Gl���c��y=O`�n�&{۲;2����ZKg� �q���a�,!_�Cg@�E3Y����DskD�ƿI���0Ԕ��đ��bd�u�/�%>n�$U�^�^���)~2m��xwJ4�<,���d���*�p�b}��%�s�:���PC`T��H>�)s���9�v��l��ӢBM JJ��_V}��4�Q;Ĺ������FNn���?ů	](��R2�[�Pe�����g����g�8�����p��~���g��]�EY����iR�=��xbǲ�5<���P�FεX&)�o�RA�/#*Q�K��~�vSDJ��;�;֒��+��[�vdy��S�<�0�g�{�aܛ|F��׵�ӣ�tp*�q�4K�_�`+:b��˲:�)�s�1�SZ1��f���|�y÷���-\u�#{�n�F?\v�����e�C)����6��>J����Hn]�F�v�̌����*��������?'r��0ŖM-��R;�˯VČE��,��:o�5��H�ä́�ͭ����&������k'���X���h��f&.%���)����켼�Q�L}�QnG�9A}
Dj�p@/'�5��E��	�˼��/�Â���ﻀ�4V͉������̦�QVH�FO����u�Q{S����W%���X�� �:^����*`��\��ޚa}f�;avb[_C>���=|�N��e����/�d�@�Z��R% �8�a��/����݇G�ýK�G7�<A�H%\'wNu��%cGEɻ"�m�V��`!����a� �����81Z�|����0T쏉Δ�e e��u�Нh�K�����A�̌E��PQ��A
S.&x4�ġa�{���Uъ���5���X1�y�f�@��?������܆lQgG�0���؜S�!��ڱc�~���2I����a��S��R������UH:��Wɺ:��BY��;]r����
� <c]j�,>}�3��oDR�zϛ�VB�2�\��Lh�K!����cr3�{b�͝Ƃ�%���"�vj��$����V���e����X��}�q����/0�� ���Xi�~�_ݙ��>bATߜN� ��*b1 ���$ �Pf��۩��DR	+/������c(���~3�,��?!+������Ÿ��>+�Ml�],�)�c����9�1�x�b�)�,V��'�}*u[���A�|<"n��Daa\����.81�O"xY�V���4�`N���`>20P,=��a��]��㺍	��QLC��@�X̡!�_�ź_�k��v+x��t�)�8�\�ɺ̼p3�ЌJOs;+9P�"-	�E�Akst��Uc�>V����7�����8Ғ��io�q|л��"�7l8�!K~'V�̇�NSm ���<�6;g��a�2��=���������9�s�sN��~�3�y D��e��=��S�����ꍩ�����VmZ^zc�R��S6o����T�/WB��t����э�6�; B6	@��~#�z������B(��v��!���R,��� ��qC3,@b*�'���4r��.���1¢m�j��Yn8w�̨�8�g�=4����-��DEX��=�ɪ=|:��T�kD������t�������uͬ#�3����vY�/�LBY�U����J<�o��?��`�m�74�TR�-(��'y��5���Z�`���i�K���}ܾ�#8	���3��@MwV:�Í���O]�*!��UC��fג��`�ϫ��B����B �Bt�(�x�feЫ�8A�g���[�l����M�p�i:��ϼ�
z�@�/S��;>�+���/�XA��e�ռ�� .��#[ɨE�[�60g:	�©QX�l)Ʋʚ�ޭ�x��&����Ǆcp"����+�ۦ���M����,�E������P�`��rV�Q�}�h,y�%��.JӳF�v�R����u��5��Jq\¡i�1>߻^���2�����Y͖_�{�̕M�C�ea�C��J"�`j5BjFP�Ϋ�M�(�0����ma��g��8&��<����eS�
8�^6��$	�CRXK�	�X�Di��t�%�[lN�}7�.�}!�tab���H˫ܘW􁱔_UNm�o�%�3�t]�I�ք9������r�+�~�-1���\��_�U�oRP�2��-�|@j�=�|���[�&2C6�f�H{~ l��������5���x�7J�f�Z��1|<�Oّ5уkA@~��ݏN!e]-��#���߂D4��h�oΗ�U��c��_�:�a)a�2�\pe1*�l:}�NZ��r�G�=C�O�l@Ax���̧]=U���>�]�hI
�L���
��O�~�b�
���	�J����>��1�Ͱ4��3��d�{��/�h�W{02Нxg��,��!y+��W�NL��̈�ª��I)��x4��*�ม*@-Px�a,��Z�����b��ķN�?p��m`Z�����9�U����o���/��S�/n��ɢ�~�D��=�x$� ��?A�	d'��d��	��~�ӡ�YoC��e��~�@S0�t�p܊�S�����CE:��A��d�M����w�-��pa������@ʒ깟Y�C��ĦB
���ڌ$Xޑ�jUz�z�n��b-/c��s�:�?`8Fu���}W���qDV�i��ԝP�W��ЃH�D
���zɱ
ВZ	�?���ʀٮhN�I�����MP,@�a�ZF\.P�`�w��hz� ���f'k�ڂ%�9:�=Գ��2>����#�h��Ű���D�f���i�}��pf�+~{B�Y2ӂ��}i�kc���	�7E�	aB�7���pYT��M%z��ñf��u9�R�)Ǻ��8f�a����[����r
Ӄ�9M�Y�CI�^�ή����� �=�O�����,MΆs�(��>���{��_����0��H�J�$�Z��E���ڿ��%�Z>�4�6壋Y^��� p���c�7���	ü��*�t����c��<1��WEO�N���{ʣ���d^,�f��w�p0�d�r�sؠB-�o���kwV��/yu1�4)�Fz��i,�v���"�`��)xf���9֯̽�
������{����E^��s�%�5�~Pv|I��1�����]>Q��[���_�<�=���NETC�#\�L�D����ɲ!�Eޘs�L�L����(a\����x4��%������yv��r�S�������mg�C޾�x"��
,HS�Ya�[=���̭o�FVt�q����O�xK�1��^�J0ق����٪3�f�����!<?f�Q���HRT��&>̆<�eRI��P�>*Kr����HĬ/���H_��?����9f�,�-���=�#�Jl�Q�0C��8
*�W��s�H%��%��f�����X�\;���>pc �p����I�5TB�n�_�y �+�s�o�,ݘ�l��BG��9��*�S��'#��HnGeg5|O�P���Ĕ��d�����Eö/ʡ��W��D�ѷ�#~)Z�"�OW@��k��Z���T ��@����1U\�J[�X���"P6�Z���2��+�;d���T��t�_��2F���ӷ���� ��r���,�=v.X������,�H��-Ã��T���A�Χ�J�äJ�dNE��)��\�㌓o�G�(i�%Xǩ�:����m������<jz�ѣh��;�sAp5'~�-���v�?	��A'i���nL�_��&�0�*�m�������[Q��X��.N?LE4�Ȣ�ף�N�\�A������D@]�BЖ&��K�e�˞��p5%,��Q���/,�~�Vr�,�r겉A
F����]��C��>�*�3�ڴh�(ql�,չ� {zjg���M��\��wY�i�W3Cl�qih�2� Lڔ�ē	�`���I_�3nd����'zA��?x���Byo�`�4�9��}0o�yiA�:w�2��k������D��|����d����wf�d @�Qt^�p�s֭��z͝�n�D��a�@��g��b,�+��wXPц�q�^�	@j�;��J4��mc4�,��1*�]ϐ�?mm��T]�����0�L�)r�=���7�_@�*�_��<��9�O�����:���ݩ]�Y9LN�
SY]Arw����zj������|M(p< ���j-�&\�ɋ�O6�	�:�!�Q��;�~�?@�#+G("t��U=����J�8�HQ���5y&�	�4r}�����D��Cn����_�2ƴB��qZ��m��?�0�?�f��.�l(�"�yz�T軇=ڐ���Q-����
��&�V)?�L|�t�`�����g*H������v�ѷ�Z#��{'5k�~�RY����k�X��9���PH�C&����9JoP���{�Ւݯ�$,T�Vؚ1*����"��Q��
�@�ܒ�ع�����uϨ�N��l���J����Y7Z�,g�콜� Ԏh��qv�����<%�>�ʐE7�Ç�+@�v�5��NH�b�-����g�I��{)͠�֞iA��A��oF%m��y@��i����Ԅ:e��+,d�P�܏yF��9�ƣ!���m-)���=D }�Dh��@����p� �[މ
�(�ֶhz<��gR	�jE����i헐�i\����V�{�k�����iXg�gqˁ�~��cU?��	��3�0V�3�;�|���\�g�'щ�Y-]6b�����_͝���ʴB�S�Q>�M,�1��}���!V���Jn�=��U=��cv���N::�8�!��qPA�s�Qڹq~����w^~�r\�vd���gC9��f�h��K���ǚ;q�)��m���2C���^�"��c����bc4����ٷ�?<�y�� �bu��DI��|X�U(��=��vd�r�T~���j4��h����*H�h`_v�9��T0��Q��:�!�v���\R�fދ��A��UaF\�4�@
������	B��B��J�)����J�6+^v�nLy�ˇ/ӳPf1F�t!��8�^˛��=�R����~7�?f��[uzn����zi3(w� �:oʭ�0���ᕹ��w�z_	� ��8M��J|)�]C��L���"�Ks���2�����E����P��T�t�&W�Cu��Y�%f����@����ۅ*o/i�&QE�TS��5i#��Z����P(���'�i�~�y��w?�լ��a�\79i4>5�`pal����X�v�'�g���_{���3f&J��g�ULVƀۑ�jޱ/��EBb�Y�LFZ����ټf�/8($-���L�1e�%4����Xt�|V�%�q�ѿ>��ݺr}�v�@FyK�}�iftޑj�ʦҖD6;n�ݺ���É�ct��� e�r�����W��ytLdh�4
K%������p\e�^f�|.���CjL{�_�q�����Y�����Ly��R8r]�0q������*x_��z~3Bh|�3��iK0%$�J��u/�i�r�NCV錰���eb�A�I�l1���Ӌ�GTO�e1Z���Tov�2!�Ғ"�~؀1�
�Xl�J�^�(��fqT������d	��K����E<�7�0O�aU�ܷ� �Z$�a�1�Jn��+��H��ɟψ�\���� ���;Ba;Q�-�m؏��4`����:��N�Z ��E�$'����� ����\{.�S���'�����Y��U<ʱ�ܯTr��uv��5�0��I�ڶ��6��Z���PApvcvt/i�+4��X�w�|m��1�|�isp��\��6�?�y׉T69�F�E�����u�>�����)�ɓ�,�&�]��Bk�����ۖ��F
�æI&�̝�k:����H�{�n���g�̒9wVF�43�D��B���)��?�$E�'��vuSo���Em���3�Z��ν�f %j�	8�|ᨨI�Q�#5�Cb��:q��|A�c�
�׺:qi�|��3n1�.ʭh�5���ڊ����ׄ`<q$���U�D}	�D�3�@q�F{х�p
���'��H���)����x0�<:��`�9;��q�YY��|�J�7��hi�׋ce">ɡ�K�SE�Fxj����Ϛ�b�u�7��u��I�K���9�M��sg{_�k��� �D�5K3���	 ����M��_��z��r�1a�b<��%"��8�}���b�a/�������I8�צ�}8�Z,���q���v���"�T�T'��"����/��L���bF�� "$.b�&��7ι��"�`�"^��LYJ�2�vLN�O��� p�(>�3 ����3�]�{��&���e���䔉�a¬�~�̺_e�ǲ�.�W�PƯ�o-��,�s��!)��դ�'ב�5�= �����0@����%����{1�E�FOa!ݩ�M����k�|	'yW�wyh�����B�[YalY�<��-���	�;F��&n	��0�:63��h�F���%�V����G���	�Y%g��*<6#=��3��������R����v�bb9X�іEUki(�C�� U���Q��fQ����ׂ�M�G���5�1��%7Ŕ��C[m�ڹ>��e"��	�����Ж�Ab�4'o���L�S���C��P�^D�%�X��۞4�J����,i��A�շf�y�t0�;5����<��nwQ!Z����m֏�Dtb����Q,�~5���N��^Ӓ�\5ogO<���;���:d�qGKʄ`X6�0B�,���&�!��잸�����X�*�T���$'�@�y#J��mϛ�|O��GI5:�L��[F,����{�	v��#u�W˄9',O��:��[�Є�;h��ۼ�5�|�;�Zm�ϐZ�{����^k���]��:f�&6���2�Z4���rQ�~�����j�*�"�_M8���7/"�|��P,�y{+�l��	P�&��N��P��|�\�>��3�����玽�H!���:��9r_""��FdD���k�8��v_���DR��-E�EQ@��K�4�^��:�EJ���''�Q���	�5�Fg9��q�b�$' OAhW�``ë�s�P 3���!}~bJ�,2a���7Ӝ��{�;jo��oW6PR|M�ޤ`o0����E�[����b�X��C�Z�N�}J�5��N�A��h�0T��o�#6gE����=i_"��4��n�]��ߡ��������M�C�d׊���ŋh L�2���s�xMŅ���:��7y�����8f2�#�y�3%��	�[�������獑)��i(�Duܓ4�<yl7!w�S�q_(����V���~��*�j�u�KG��j_��A T��w��[�
��G��z�q�-v�g��*���w�����T��r�'�(I*T�!2�Τp���~ xW�"~�W7�~+ߘ	�p��de��9�'���ե���շ�CTR�Ў���l:���i1Ǎ͠3:�8k8ѝVF�&��ѳ*x��9��m��k�N�v�0ڛ�����P1�L���<H8�;�#K�%�D%�*x���?��2 ���j�~�m�r�K�-4R]:P�<;��
}s(����T�M�2/�7�?��g��q�z�:Щ��F��\�Ӟ��`b�0Q��Ca2���2�;˥���݃�c�K$]<�M�1��F��N��TLQ!��W�jZT �Q翎rLx����]�eղEIF�����3����������K�-�s�}���V����(`cj�@��C����j��W�1�[Uc&8�u��.���\�E�5�2�X��pc�+�����P��7�a
���`��x��S�`�շ�M����uU�&W���ŉ�e���&�MW~�@�;���ɔ���Px��]TH�����|x[�FEO�*,���}r
�\�_�]��Ȏη�"���~
v����ׇ6-�]dK���Q���O�)�8��n���n=%�[�R;*�A�����^ӧ*!)�[�F'ɣ��R��8!�6���~O���x��BM\4L�B�N$��9����oca�㮘��:߬��F�����=�K*3ie8I��5��,�0xR���J�(�� Pe+�7���1�����w�E�`�Lcx\�F=�ˤ%��j���D��12�Q����.�h��8��<ѳ��(�]��cn(a	U����9�0��$u�ba�̫ڍNBu���y�Q���
K���%�c�J�[�7�󽜛�V�9��� ����P33�t��Ut|�H?�+$�XQ���#v%(Ѻ�Qm��po�1��X��c�Yh�|\fy�V�]�$��E� ���+��F$9�|�*E �9����M���ώ�Vx���򸨞���M&���MX�F�1����y���њ&�;��K*ٔs�b�{s��l��*#�F�ϥ,ux��� �N\<��ddQ�������Mӛ�b{�m��L���>����U'!g��������F�?��0�3֫E;�62�2��񞣟���!~�|�kU��Lƀ�����[k~ )#�;�F�S.M�{^~�J��v�U��W�<��{:��	T�Tf�/��O:�w^�������Õ������Ov\�F*��N�v>�QL�Y�"���@)7I�\@��=��vW�2$� 2;��Ok@�ț�h�_N6�ST0�5�n����f�i]�w�X�v��m������"��֊��C��TOy�m�
�ӝM��*Xi���v'�{[la8���6H�2��ߊ����d>Y
�@}0W�ς�1
�rY�|��i5�_�vB>Z���V�\0���U�`%|�0�S��s˙�:GԪs�@���.��� �*���t�܂��	
R�F�@m�5C�����4oA�C����H�Ra�@���9)����d�loH�n��@IB��t�)��ЕNl�-�X�Ƥ�S:'����ۮvO6I�}��{Ʊ٥s�衠]@L��b\UG�ĽBmL6���p��G���f�B�ǎ$��|�Vˀ%���!��3/�p��3]:O�28��
��y��P>�J��V�J^���Ēs��Ɍ��y?����6�u}�PR�*�2y9^]<Vx�C+�P��fK5f�Xq�ʙ�Ԥ�v����r�y;q��[���Jd��~���g�����U�Ymգ7E6(mνYi�����eenhX��1�gw6W~��հYnY�'ER��>E�A�������fs���V���<K�&[�<�������Ym�.,��P4��E�X�h���s����E��FH1�btq3{�{�Jc���P#4��R���B�T9�����݌$���ܖ��Cǉ5�y��a������-���Z���5]��
u��.˩���#�:!-@��](n|��c�A�h,C�s��nf1;�J~4�8��당�S�I�k�E<����d�d��|�G9BXp�r��\�h:��� ��!JE�sL�X��.��w\����JS�Q'����cVY�{�)&p�bM�iM��3sa����8�d��w����Z��'��%u���{9:�I����+Te�g��K�T"c�e���m��#r�so�FV?J��U.���`8��S�1 \9���
�Ʉ�.VK���z�Wt�)�T6$�>��) xyi�>UP.��!E\�I2M<�MF�1m-'h��w��Uӡ���9�Ն-[�Ɲb�J�L��y�hꘖ��q���>�����|�.nE�1g׊�$4iM�k3���ݩ[KR��ou�D&#߳�'[�M�*��4��ڹ�M�K\��u�4w	x�q�� p�+%qy���π�H~�CJ��X�0�q-X�X�N�f����Hb��\�Y�b0k��Y�ۄVH��][���僜W�AA6���ǵ����7y��������x�5�6�icǧ'��K	C�0葏�D�G�Z��+��E9��i�h�' j�4)r���"B���F�!�Л�!AGz?��Nt�K0�P��U�	��i9i��) �cc�`��~�*�O�W������M���#�"���o�@jgmn�TC�%��=g�c�����!�y�`�iWg�s�$!9g�8�d��o�l� ��h裧WԼ>g�����T@�j�+ J2�K��~���^�a��wBP%)ys����2�7��u�E�l^���!Aa���v����#|4��B��s7�q��2x�K�J��
b3Sj6��i�u�M<!!�����0Rg����'\��#s�Ŗ�eZ����a6O��я�G��W�H�����`���� �OR��4��:������c�߰�@OǙ�|V+N����\U�7J��T2`s� 6�-�v1��d_&뜆=���b�&;HO����)�?^v�"I2��B�.Џ.�K�����?��.��y��ҁx2���%�it�t�8%��L��<���{)�;���C���3Z(=�rJ||y��)����%|�eD,K����g\����r��W�|��v�)Fm̓��0PO]�%�=��iaz�E:r�b��-�2z�'PQ8�ǿ��ZUp�y�Zݛ]?�Dg[D�NK~u�>�����w�/���}������v|��xT�ԥ3���X��PR�� ���n�%�����DX�b�L���@��~���U<����ҷ%���V�m�'EA�)�"-���,�-2n3�M�."Ð>�� �Tɽ�I�P�Γ��4��|S�, �)��0�����G��7=V�e\�ԡ�{�?����7р��00�m�r�r�b� ���qU6u�s���@-b�4��#�����5�Wgd4�P��;㻿|�#���?����4X��<kC�JGEм��u{�?��t��7����H&+c�hEUi�%O:r�g��%�[ñ�O�f9����Ia�Ho������Rc]�@���SU�V	��-�s8@�ċTvwe���E���a53��W{�N�D��V��:�g[ �g>2��n��]��R�mY��b���ocK �@�ǎ�QX���i�g8{7ȅG<�#�@ᑎ�@�B�`��"ǉ�ugm�))�6���E��ՠ�J�E��������z4W���(���s/j$+0��9L4�y1t��X���
���[t���փ��Z�kA�F

R�~��%�ª�s!��uqb������ܗ��b/'��;G�1x.�������,b������y<W�'�(�T3���␧�����oM�m�1��X�ۤdQ���<�^&�]߯ �z�/b����?�ٕ!�48���w;!1���Cc�H �=f�e��f�'�y*�;3�ѫ0(��G��X��Z�-��u������疵]m,�,������t���q�l��BT�<c�z~a���E<�CA+��ku!�|�0���0z�ЋW�hKZ��� �4%gs�||��h��1�#<�'������&�l��ݛ����x�F�;�	pgՊ��.'e�>c`s� �[Ljܻ��E(��n|��MҌ������8Z������V�3�"�����{��tў��f�efvvo`�^��K����W|��$j��ku,؉��"�%i��J̳J,!���&��0?{�0R��cxbq�>�B���v�:���R=JI�}�����8t�g�0��
G&.I�2�������:��_��h ���$���E�-�Z\��	�f�<���D��� zK��,A������dZ�Ą ��m���
���i��,؛^*���hЮMϬ��� ��?���ɭ�Zv:׊�Rm��Re+�Cn��V?,Fŏ��Ӂ(|��&A)I�N& ��Ϲ�U�Ia�����}���g,�,�2��6�{2���|����!�����_��6�)��[@�?B3�I׉A�ߔ9?D\�җ*�sfa�h�`O���"�� r��t�Et�����\)9��%n�d�AV|�ـ��<$/�&�,eŁ1e��|�P��^�5��E�03���p<�p� �K]������Wz�:T\O�ҺZ)���eO��o?�b�.�����M˥�C�G�p����y�?JA� �p���s]�X��h����#5��n>�z�i�k8�:�e֠Ĝ
�1kx~O�%� �%-)�Ea�U?_Ĳ��&��_����x2�n��\�ɬG��~�nT[�
ɢR25��òߺV��@��畾���,��9832mi2Fj�iB����&&� ��j3���k�uC'vԠ�"�R.�8/�ФqX�W�o�5k��մ�������Y�F�E�4FhQ�v2z8�B�5�IN�_�ҿ��W�䍟�l��f�ą�Ѵ+V���D�C��7�O�D��o�p�:��3*����� x���<v{��4�B7�'Me"!q���-��=O��Kps���X�����[�6�Rs����c.\U��ol� �59֖{�5N��0��MI�<�]{d{2�l�L��1E�K�A$}Aޑx�i��ݦ����#(��o��Rٌ�(�3e�]\��9�dᘷ}[���|KY%������"gШ���iaNe��}�7���̇�d�cg��Gqz-���cb�����2X���S����{>ؠ��:�.�A9�$�q�M�ن ��\ ��7�`=3�{�'��W�1��ަـ�˲����Ȕ��ϗ8H+�8�3\cJ�y�tƆ�����>*��KW"]4���p&3�k�(�k�-��M�����)��v��eRR�Aَ�AŦ�D�\%t�m���$�����Nx���u�'q�am ������JA���n��X�\M��( oЁC^.â�g�=1�Xs���(��|t����e�|��v��()�OX/s�AP��&�9���E�Ҡ�0ʌ;Te��nt�t��nJg�ea�	EP?�i(	u��W�q�]��㡁c��dz����P;�?�^6���}`�vW�~i���gۧ�N�	�ܦ�ˏ���� �V�L�#� փ����^((C��3�a4\�,t(G׶���$�_t�O��9�mmn7U�9�5#t�% k]f���޳{�_I�MHY,h0���V����~�^>%u�C�D��x��p�b/@P/F/�Tm5����bU1���P�R��|�('�N��3L�.L���x"D��C9����v���+c7W��1Ͷ�����F��[�[y{,5c[��,ȿ��d���.vi�`�f�b�\�(�L���YH��CCYy'2l��5�#��}+�"����ۅ�_��֖��I�VT���l�o��oӴxd��E�m�c��>6w��
p����mO����¸g�z�����<��W�Pq#�*�m�~����#>�|Ԓ�[3��w��+b��q�qB(�L
W'���1�Y=����x�]�4j�*JH����JT%��[��SV:h'�CB�]�d8 8 x`4v�s`�c:q��ٖ�N+���$�K|	��!q�,�2�F&�\����:���۶(V�0�/{�ed��f��G����d$Xۂd)�r1R�I��g���u��ψ���Ӡ���iH��E+�IC�К}����]��夿�+�7o$=��~I�%shs[�d`I�{�mB?�$AO�U)(
,�G`.b�ҭNb�j����� �@<4�����S�� ��̄�T͚SP8��{Oo>U|�7��=pi��:������N���k��;·�~I�s��Ts�&~.!8�j���jZ�Φr_4�o�d�D��NDj«�C�jH�d����x�QBqN���յ��������Yv5O�=��e��'��0�$�Rￄ0�xp�0��H#�<*I�9;%�Y�E��	.���22ij�A����Gi��`ms����:;���#jN�'^q���3���g��Ś�i��T�/�����%��(;�-��<"�"�_�Bý�a�4�D9������j&߹U�8��ٴ�F)zY�?i@`���U)������h�!Ґ�Q���r����b����8nq�/ppP��;%��G�W��Q�[5Vc�'�FI/��H��y�(�a��㙙�򢨳R��
�C�ֲ�\�;�bh
�iK�� Lf���@�����������h	��ۛm~`�)�ww1(2�d$��/o�����8e��Bc���Kb9�Y�+Q|���&������QRL]|X���4�OH���1�<���-e�������4�ȳL#v6�$��bR���gJf��d0b�|�'cj��k�ÿ��ڨ���F
�(i4�ր��44p����S��}���	F��Z����|�r��gO��浀�1މ�/��S�q�<���o[/ Zȹ��r?��V�ԛoU�-Pє��/}k��Q%�C[(T��M	�L����4
�F��$��|qf����Y�������}���g��Rl�����JC0�a�΁��.��ʊ�hVLrm���ݞF7��@��6��&mM�ܰ�O��A���}���[n�R�!k��-�0B�^�@�G��c�~��o�N��G��~�cp��L��I�"ע�6EK'E����O�攎���r���c��i_R ��A�>@��=�DIw��o5��"�ѵ���t.�P%�e�J����-J�G����5�%y&�z/���*	�_B+4��'N�k��|� &��N�9)���[�>:gq�
!d�[Or\��(����6�c*	�e���&
3��~2*�
��ݏ��&����ۼ%g֤~�/q�cdW�+ŝB�r)�?xrb÷���D��=��R_�&��e�Gˠ��8bN����!��g��Y$3̆]�m�כ����,ei�(gx�#�OQ����3�2A�	4
���q����\2.��-�N��d��-����د�ɨRb{M�1r�b���鈇��Px,?~M��C*g���rҁ��o�����r.����8)q�q,���U'�3��?a�����b�R��
 kn\З�"�AyI�M"����;�0r؄FraŰ�����)��K��c]�N��g�ĬKG'R�){A�$?�M���Y~����1���l5/�\w��ٞ&	.[+�~�C��F�z��i)X��ΤZ�_��ߵ�%��c�w���{����W0 ����)AC	��x1�\��d���y{֬|?�q�q޽�<蟙h�C��vݦ6��8�G�Ӥ�8��'���pU+���P�� A�^L4�xf���!>	��Ք����B�~oͱ���ϕS1Ht���9>Ʒ�5{�Y�#m��Zg���C�C��4�>��4�%����:���4�!�Wy��q=ϼ��j�w+$#���#_� �D4�ssU�(�X�5���e]�e�"����i�B����m���J�U���*v�fg36&��]�ۢ}����k=�Y�$=�2� u>����?�W�N1RL9F�8���2jD�����WOw&͉�8^J�l1���?|��8c�����>�v�*��k��?�J��Y������Rg(�(.,5�^�PIY�:?	"��,�����\��Z�������&�!U�t���;�2F����v-V:�g��Lo�.F5�q��Dݶ����p�3�=J��;0;t�m��ˤ�K|�A�ֵ�ĳ-�c��#U@��7�BLA݉��֑����&�՚�������u�O9m(0#"�v�����l�#����m3��,Hx�.C��D�R�]i=jڗׅ4���>D��E��
e5LI���?���nоFw�Iə�(>���h�<��_S��D��G.�O�տ�-��	�
��՝@j���G7��0�x�V�}ZA�2�.��6h�]�R`��%3�@�Lk����6fѿ�Z�x�	��r�U���檦�BEk�/Zs%��~��w����@��Nh`���"�K�'2+�	�\���5-12�=�6f���N�<T�aj��O��]Fq��0�Ll�Gܤ�tLTX����r��q"�<�����"`�9���}�ɑ^��x{�lVLC�$n�~2�-y��+A /��3�!F�se������p�0��m��a�?R-;�ź����`�x�w��Pk'ͧ4|`H�;��f�*�@�CV��EN,}��}ە�M�3h�g���H��ҋ/
%pn�8?|I)���L�>�#Ma�wd�x�*�j\ݤ(�?8Q��q\}��䤫��j躒@��)�~"Ĳ�9�Y���y�$��XP�E$���Rɴ�7O��Y8EPǶ����/�����	�)�/�`��G@��}a��J�y46�콪W��k��uN8��I�Hc�c�Z���( NP�R��{�m�AA_�T(���+��p���*h�߼oLc��#��[�,��!�յ�4�\��Y�
"�F���B��m25X��֔����|�>?����bߘ ���W.Kru�a3U��v�1��y�:��x����A�%���!���\	��XV�,sӭr;��q�l7dp�`AN�Ѐ}���_��D=����9���Y;�m=���$҃z�c��ꆜ0��D[i�tO0�F�P`r$`D�b�څ]��?'ѹ@9�g�N�A^)��1� x[�3�HP������ԚQ̿�?ݸl�L�@9�/a���G��)��2VT/��Fjs���`�BLW���j�T0Ӏ�f��#����93���*&��	����7�1B�D�(��=<A����iC�J0�;�V,�J��kO*9zE��BVD���o��#E�O|�X5��Uh�Ha�>U ��ἃ��#�%��Đ2�p�E��F�G �a~�N�{���0k�1"뮞�̆�F�:C|��j<Ώ<~ ��:.R�}H�~�&����
�߈��R���B�q�	��en�z��b���F����M�]��ˎ|z�2%�X9�!{>0E\V���D�!=�ￂ�ֿnx���z B)�z�OD-�� Fis�)'2�)\�}%s�����&%��g���nD�4J��Z �D��*�5��X��ŸB�pT<zb�)*��WLŬm�����Y�s;�J����t�����j:�K���?Ҫ�d��7<�
O�ok'�q���1g�{s��Y���.aD�^���&�����9ҽ��	v���_Yt2���qd���$.�~#���
����	������(n��C!��[��D�'��J�+��G{!��G�˭��S�!.�<eŌ�5D`�ʮ��r&��P�I�R���߁%��`;�M���-����H��8�EM^
ocQ���O����J�r����[2���؞I�� "�@��,-�&i��60Tq\g��~g����З�`j��%�{N��决<#�5H}j���k��n�EZ�u[��	T�%ȼ���M��0I=�`K�#:v�S���C��/��M��r�@T�ɀ�m���ȯ��=P�$}�K�DM�R���&p�?��"J�[�~Sh �Ǔ�D�}$
3fx�n�u��P��!K�E��b�����Q�_��H��0S�~���S�L%��_5jK3�s%�J���P\�X2$�,��RI�C�����k�7�����nc���VX���7�����rX���a����pڿ����m$~0��@��D/�~S{J��1�%�s�Ŭ�"���ם�a~�|����B)���?'T86G��I]���(峮n����$�K����a[���p57@ߚ39*!���Ek��E�~h��8P��U�� ��ǧ�6~N�>��fF㰭UDe2\�h?t��$�w�<���n�$3�H�5��-Ի�"�G`�n�l�뺖ip}�a�HI﬊�����?|�� e��aF�d��K��E��}r�4w�ߤ���(g����1�󏌂�x<UHCb����s;?����7���ȡ�̏O��]��5=��x��}���4�����Y���6ՏQ"yb�I���\�� �t��lq.{�@��@��%x+���MaT!�:�C����՟cX�L��E�\�G��MӠc���W���@=�욌�͐�Rv��_kf�mC�����Q?�[�F`���^M�W?W����,�]N�ܻoCr(��Wɔ�N��f�1�Ti�	.�鹕�3.ǋlP��1{�ֿ������C`���avOnm:!^հRi�3�f9'?.�b�;���+i�j�:�JҾ���ݻ���xP=s�V�Y�AHe1�O��$��U������Y��� �Pccczl�w�6���ty�93M���Ɣ�2�4��I-���َZ��,�ѝU��)�q��8<��k�L���g.�(h���1n'~�K���sc�(h�y��<�&���?�K��+�hS�?=�z�'l�Ν���ju�G������<Z7��(AT!��ۘ�M��6��PS�g#v��t=�:�gU�a��p��(�������i�?�ɕ�����cK����?Oz ��E��H��4n;��R�x�mcrh���׻��++"�A�����t���Z��T �G�J �ȓ)r����q:�6�����;�a����K�B%�ej�Oe�!���hT�/2�y[rHȸ���[�yJ�g��)���NN�E�h+[3�@[��>L��(���D�J�|�O� ?&�#|��]��/���!�;Q���t�-[@~ ����P{��R[��Q� ^i��`(~�ݹ��7�ݻ%�yi�ԞQ4��xO�`l��2�atY�:jV�@�t�N%E�Q�A�/��w�l������>�V�y�<����j��:�v���K��'e���W�<<�ZO�Ni��ܟCe;�� A�?�K��dQ?̐�V�	h�:
������B��Y2j8���k?��$2��\���W��w��w���̊�|�)^8��g�i=�02I����
k�+��}�{��u����K��`g\`��+l�=>��1���\d��F38h|oi^T��C>P���v�!5ЊH�+Erb�+�^��-z?N���3"/��?��py�dzp?h���3�D�0�t7��Ͽ���m�w�y��c:}�AT��N$��'b���0����*-���w�� �軟:��U	*x�\�1� �ƒ�̦�-v�lv�h��_7sL)z:/�+x���0����I�W�cd�uIŊ�J�>��D�����y9ˉ�MQA�t��@?��w��P��q�ai`�6ěw1�{���K���?�}u����Q�c i�ͅ�z���	�J�5����rŇ���~p�-$��C�Y`*�^��/ܖw\�ux0�B���.�,��0 �Bŀ��F���iLB���~)��L�1��U�YY�3H̤���0�g�@���\o��O�ܐ�g��6�]��� [\�TEL��m:��T.���+��fu^5q���4���{��C�d:��E0nz�I'�|l�(���q ���3�b1k!V�H��:�(:��ޙ�d9���J���?_�����qC-�;�VUzˏ��JS����g�-�b�a�]_A�V�C����쨁hK��J�n�6����̭Ed\T�~�O "�����*�bRC����U��đ���W�;�������(#��d��y��잛�Z::�20�/
����r���]��~��{MFL�}Sn�D�k^MΤJ��:	e�/boY55��mڎ��	�]�t��S�j�)p����~P&�����w��y��w�l�g��$�Z%5j��frqxI뾈a��lq����P�4+�Z��'1/<�|�F`��gm�.�°gd磏[�2�/r$�|�j���_�[$P���pd �0�`�I��	A�i��kgx�Z��4F\1g+��
�����]���"�V�X�� ��|�	3�rR�_r�Y2e�����d��'�4���a��|N�P�	&���P���Gm�eqX�#�YDsq���b�m��[���b��O�����~S��$�����.c�&�~��U��v^�r[H\��y�>�����@~��h�[��O-�}��P%7j���lh���J�NBR�j�A�~���,�k��^k��M˷&מS�N]�ئ��#�ڜ�}~�'�����T"�
h֜�N��<���F�*7�B!d��!5�v�x��ӈMN\����A�u͗l����.�:8��(��5����2:Aá��Q�h��fXk@��O=�"��R\}������yF $[�N��5f��ӌ�᱀�VO�$Vc����N~ǒ��"2��U�g�����Z�.���".$k?H"���f5-�.}�EW���-��j�_V9��.��e�F�̝Ϥ��7Op!�y.�ȵ���Hb0G	� �L��2:���+�lX��C�{I[��3KN��j�T�<�U���
~m��.3q�����;2�a��ԕ���[�]u�$�2�������46*qH|8L_��ީ�X��eh�Z�&��QĂ�rOĂ0��2y+qsb���N�)�P�QO�q�i�Ч �&�,|+�}�~�ԁ��X�����:�!/T둀���u�H���a����Ì=��C�|Zv> �^y�iY����9�%/ ��ݨ�P���jY&����ђ�}���'���ܶ�!��ѽVc����g�ݤ 8U�]�J���+�B��)�h�p#И�FHQ=
NK����4A5�]jp�.2��n�������8��I�V�Y�����2xO��(���{���ęBt��ln©Tk��CK�vف�Q4��Ը�-sj���f�㖺�䤀�5V囮��n�]�����r<�,7�od������M��K4!dZ��U�e�&_����v�M�m�>�+5 )p
���(=�����Q�V_8u,��j��'��]�b:kMrb�i�B<lM��G'���~~��C��>�@����W�ӵ�K���%�,����W��oQ�A�lV�D�6�&P�uM@���	�"@yZ�E���FL���4�5��e;\H�!������>�<sQ}�E"^G�Q�U�/���5��q����yv����p1�'`����NꂧN�&cz.�)���wɊ/佈�9�N��_���U�+�qD�4H!3��t�*���K�	e�����G���Bð�Ϫ�H��w�!��3��,����^�O(�]�J��>�d��ڂ���@�la�v&��b��Us��neߗ�4s�»K$�ޗ��"����<�2Q�M����U�)�J "���@���.E�S0�s���A��|弧�+�Q�,t÷�Id|{�z��~O�����U��Rw���a�=��W8q�
K�N��GX�?����`z�v��1%6Â�*�I��0ךt��N�����O��_�9Z�X���ga�࿡��.�F���fO�T�sI�����תѕ=pQ�];UM��/h��[�~l��%^��t4��!��:��l%>`�-{��jU��<p\}�
�ǯ��w,����xb�g����_�_��%�$L�چ|m恮���y������w�*w�YY�qn� ��������,��}J
l����'y�q��0?������{����vΔ��������G�J��fAj6��)����0u���E�c���E�J��~n�A����(��V0� 
ɜ4
utr}�����œQ *�	�r�$���;R��o<"�h�S���d��ؽ��_�{Ҳ<]A�9v�U�ɋP���(�Q"�O<x�1})}8���cN[vO�!]o����4�/ [H��]y�}�h�n]-@�����ԫR��)��,6���m�0�߼j��Ԁi�qͅ�P����f�&
�5��*���k�9�����F�;��>��l,�:��3��� C��8��Q�\����]"� �k.ٖlV����S/0��7JX?��U�[5[@x��޳���}�]�����qfI�t�4;�ѐ���"�C� ��x��h+n'*�k�4 �E�ͩ����zJ;�%��b���K�
J�{h�[���ıX�5t��ȃ�lr�7�!js���hX��zGN|F��f�[����0�,�ٲv?v==Sֽ�v��Q�#�NJ��T�����Qa��x�O!��/p~�
Bm�
3�t�ڳd/r�+�X5"��JQ-%2��#����v}������WnM˨N�t��mmM��D[ �We` A=~Wϗ�����l�\u+.R��Aig���:�׾"?/jU&[��`���7��=�+s��\(�fW��bF�ò�N�B��R��?ٙ��H�.���FC�=���������Q�MGUMR����׮��fS�w�y'B?��G̔,?�����*��&�ѹ4i|}-�P_v�Mp
7��g�uj̓y|N���� �h��"��-��E�a���ce��X\��Q~%9W&��o��7)�^���(�D��yl������\Sz��3[Ạ��<�c�k�π�f.mʪ�l����TN�7i�w߂-V�s�B�`�b2.X�6�uI��@�����*�珅��E���0#�Rx���;�"�t�����7�w�6�9+���ٳ�& j����L�?MOt�P�����:A������6�����T.�@��V&�3{+n�=|�*&�����\��P��xQ��	��k�1���u���V���i�k�pSh\�~B�
K7y�R��fxI�F��B�Z�>L�����
xׁ�K�WD���ǲ*���X�_�m�hL�Z@�v�f���&�HR�P똜">lk���1�,�lt���	.����xN��h���LT�����#$�S�|����|�v*}��I�?MD�"Dn<2�F#�h[Vڨz�K��7��kF�T5�>��&Y���B��-�+$�#/�[�3�L��S��+`O��m\1��2id���+-����G�o�-&�n�Q���TBЎ��S��J����M���s���� �
�G+� �g�W�=5pa�?z�����p�J��C�P�ӿx���M�W��2Avpp[y]��4Ld��Q�l�}n��>'UL}]���N-�����a.I�4�:"��N+���'��3�S��YW�#`I����'��&�s�(���hZ:\�&4A��P�猎���:ʛX��J��\��B/��nȒʔ���躿}%��=�U�u"�������� 9�ϛ��U�!0�]� ŵ9z:O��hyN�-i5&=�S_��8�=&����l�}������p� �	�Ɛ���$�B����Ϭ"�g�AN����<�\h�lLd�m� �$&��E
��U�q������rm&�;��9"P��?��[�<������i'Xj �	���5���`w��NS7F��+|���Z5w�#�x�˺�<�
㒒�>^�0��t@4�s��[���5v���w�v�͟c�)� 䄫�I�U�I�#ȫ�͌�*�_>�²����5'�9]p6��͢T.r��e5L( �DRȖ�$�sn���="q/���},�-=��b�F���*q{RK�8��B/;{��В}��3��~�~o�m]��;�jh$Ӗ�X�ㅰ�E!�<�&����	ȪLw��m?Zi�l�3��9�ɷ%�U�N��0�@hՔ|D���!۵)o�" ֜�5o���.
^o�Eo����S޹��������
�JAhO���:��s�v@`>W��<�o�;É�	�t��b]�4Ch9�
U1!}�߶N��z�&�o3�����9�R}l������0��q�bS� ��q�g� N-�2��=����l�3��f����nno<�(PMʬ�(��LV�l4J�x���7�����4�{� ]�Κ���㻧����(M�>���Ӱ�J��"��X���<@/����:���Ev`ܧ�Хl�Գ5��~n������Ag�������.b;��Gw$�h���O�/�)n7�Vަ��D���H�	lH����E*��j���br���s��7j��;���5"���O�S2%~sz�sBo}t�i��(�Z/�?i���u�����Z������tƦf�k!�O�p�9����4�r���0b(��N�=��ه�9���5?���l��bLK�O��6M�b�Z�m�4�Ht�TG=%����:�4Z���z��S�n0�n��ʘV�ü�)�S�}�ׄ�b��yר}����)���G�>�<JG{��#�iX�c��Ď*oHTGJ{���l���H���sެwߊ��8�,��l�U飹�E@�.6$!��w	_n1 R������5ԏ�����m`(�J�BF�D��-����ݺ
Ұr6�B����.���դ-�j&J�,����@,��ܰ���;^�y�����"Rs6�"�j+{F"-X���#�e�u,Z�Q5�r7��}��Q�#��'1_�p��5��mw��;lV�v�|ɉ�X�]�
��}��	@4Eo���F�Tg���`�D��ޢ~���B�[Z���4غB����G�)�SWHPÇx5��N�*-�=ԟV�pZ��(SCt�m��lA�Jێ��?>�Q�VSr@��}�����pZ�U���ٜ��Ix��?���ǛI[ �1�E�R4�y"0_��
j/��Ί�Ǥ�`w̸4xS����,D�<��&�`I�fy�q��!x����|=_���SYm	К�ԩ��_���	���5 �bO���	2���@��-v�ZT��9�f_��|{*�!j[�s�n����p��'�r����.u9*)?e�8	��ǳ
�"бN2��sO��ʻ���ꛛ��H/aڍ*=YWC[�0�j�d�\qR7�'ǅ�>�'��H(��Zċ����A$譻��K	0���P���KlD�� ��mбt��1�*��RЯ4�kի>�M�?�-'�h�!]�p��Ow��O�-�o��`��+-��U�n�������t�qNw���7(�A��G��/
W啱�У�uf�M{����;�wN����{�<�в8��*«|[d!N�whM�l;�̔T ����m���9;a $�2>������΂.��'�l�u�����'<�+�L��~�2�!�Z�ۤ���~���p<�ñEԎw�"��~{�QGX>�f�T>s�6+��/�zd@g���T|O���������X��+^S �e;� {�L���|.M��ҡ>��9���&Z{!9�$e�2�N�UA&^�Tl�\�6��it'��K���<�N(�8Y��K��Bh
A*�k��/�"�l�:7���嬂XQQ������~7@^� �R�S�2��/o�lS��QH�t?]��qEuT徭�[̾�2͈Q�I:ȼ�nڴ�������c���z��}:G��o��Y^ѨU2��.���>�v�媄��0�@lʲ8I��!q��]�����������AѼ�'�Y���;�߄0	D��^&O��R��te����KH[�9��?ò�w��\E)�H�5`Mt��1��-`YQݩj�GZ�U�>J��Yd�6�f`G1�'	� �FJ��G��n��6���v1�;&
Wh#G���ZG>���Nj~�)�����r<Ҿ�x�	:��"}-ƿ%:bz=K�X�Jg����xhG�a6
���-q�o��<֛�T��mf�Ly��xd�b;=j�	�U��Y�B�QȀ�����^���Sn�����J_���N�<��b��t���䠭�q<-�Ӆ�������{VT�'���F�P>�M}3�<���>%�Ŭ�2"���"; ��p��z[;���+դ�t�D�r���凸б������9���A�e��V�	ˏz�s|�|+9��}f�d�.\�(e�zwF�H��u2�RE�� ����Lޫm?��Ho�dYr��>A��2e
{.��e��}���κw��_jqc�h�E�|���q7c{��`C�~A	�o���1\�Ҿ)����I�m}��p���c�c=���<X6�8º���ꂡ#������O���9�K	����׍}� Z��GI*�"��cv�+ �~T��֕�|*`S�M�|]
QE���ͪ]�i��|��G]�.X�b5[N�t15�s�x2�~q�ym�b�B���4�
���'1�
E��:���d1�i�x��Ip1�X���M�yE�Pa�� �$7�}���ֻ��lo�r�ch�"\B�:���� ��"yz	zb�:�LX[��oLy�i7S#�����������;��4��Kj�"�<8!��N4�=F#Ť}=�m#!��GL�WV�(9�x9a8�V�%�z�����ΐ�5 �!����5������I|2�� ������>�a��Z�8�c�Qo,b4_)�+�5q쥍�ʫX�]����z,�=iSLN����kg`6��� ��N�`F��-ڻ	=��n_��PQ&��G�`��B���.�ӕ>�.�&,'����4��(vXF����@���6��W�]��>�Y�'��̍�kę��\�
Q[�j�gi�%�CF��*7u9!�3࿹BY:Bj-����G>�8L?�o�XCy�3 ?�	�`�`BT@p�܋ ��.���q�*�U�n��!�`���e$ȍ�E�"]9���cלu,�G��-��:k�/'|_]�ڰ��Oy�r�E���ř>���Z��;�\�GM��t�΃a�4mW�*�	"W3�0��������Q{4���a�mG�?]����t�I�NO姂�ӹ8���_���>�$ֹGlY�:�����;�[V$�ٿ�����87?�jo,�X�+�t��_��A�;��8DXv\��G��*��Evz�R��m�̲>��a�Ԃ$��g;z b���⢻�ء�B.�.�d���cu�f�0F�Byι
�7V'z��K��/��N5o �]:y\��8�.9���k�<&��gc<ª�@�yF��E��M� �����@M�3t��>��|N;:�������p�\��q�1��è��uGƝG!̰��+˽U�]H� �p������]o�G`m`s��\����#D����<BKk��m�C.��#�uK��B�ǌ��
mg����J�>������R�t�~�]4p�A]�&4;	|%��y�o�!�U�����/f�j�����ː�8'�M�W�N��h��A�&R���*����a�iC妪?$9u��ȓ��{o�a�����T?2Z-�*t�㩰;�Ez^?��\�����<y����8]��Ox���l��8,�Y�`pK�q�s���r��IT����q8Q'�|��� 6�D@;d߯�<eUkaj���E,����i��
o���aV�-�1�&� ��^Ҟ;���^��|^��o_	�W����U��ӗ�)ꀗ����;��x:�lu��Һ��o:.�=v칼Rf[r�,��Bq�`�<K�3jI^ �T�H0U�Y��]���<�� �p�!u>�[e�sv��|Q�^ee�	�sGӁ��qc��P����z[J��(��eaGҺH:y� �*���g��V��_���
�5W����L��%��;�����΋�RftJ�dR����tNM�g����q(��b@)�זӮ��G��u���cw���R�%���9�L$z��1��J�,��H�x��# �P3���i@����X��`��z_�EG�;��@�����ft	��C�KɐiUWN�w2�	i}�t,E;6r�{���O
B�?|�����+�'���e���]<��+�O�"m��@& ��`e󂨞m�du��J�)��]@dPA�.4�+�x{V8M�o��ڇ��bQ��@�~o��=�A��u[Ӷ���~L��
$q�*�lNC�e%�(�Mh�Þ��4���"1�߶���5�Rc����ű���k�!@�H~�w��ٴ,��9{Y�[��gN96ꌯ��SIS��J09���Z~g��H!�۵��2���yI(x�@�O�F��;�C���o����O!�<1`�w��9���E7ތ�Ip�TH��m��o�.���Tl�����;ӳ;�g��Ƀ'��b���,M��<��:o�O���ɪ��n���,eT-\�� ����-s6:<>eJ�E����ܮ;�ŭԯ|hZ����Հ3vs@z@���(Aw/�����
���?\�H�%ʪ�3�9Y6���N6�@
���s�k&�̭F�p��ޏ��u������ ���P����?jz}_�58+C)�5M�o5Hޖ��3�&G��H�sz.���k���:��h]uN	�\n#-�4���ș����_�"s��*�yy2#E?�s��3���G�ɠ4M6e��D�}���ٜ�3���e������C)1��C  �Ev{�1+�uIJ�=��&W:Я�霌��nSѧ*�&ju�&8�	�?�ƒsq)y@���8��,���D���d�����_�Z�y�����?ذs�Ԡ}����}y#�0+LK��<��nZ!����d�]��}��sO�;�3�_��Yp[��ɉ&�n�Z��A4��/��	�6B$��;����}Y��es�?�?1(��_��Tz�vIH��٭"5�m��ɶ)`H�v+Ɲc4��U���Kލ�o��cm�s43����|^��cspC�E��\¡����r;}���#V"��i�9��ׁ����#���&���E3h�#�:���9?�=2��N��W�3?=Z�f��H6գcX	�n��u	ľ�[n*�D5�ԕUr�ݻU�$��qFc�F܏���-/=hǛk4lS l��/��9\Q�lڗ{t�~ꓛ���}叼5�����<��lE�g/d��Pqm[�$-1� ����^L��#b��LCJW�����H 7^��@ )��ˏ�a��(ԲEslH9��.y����m�ׄP7��Z�H�",��mY5�<c Dث<
9�A)���-&9���� �Ö����1o�-�:�,�g����MA/jȲ7�m&,���`i,�]Rѽu��^�:]L���	��.����}����L�AST�=�0�?/�C��|e%��
��X���4E��S�%��Xs|-��S��HF�`� ��\���Wg�̢����)^�9J�~)ܜ�i����O
Z)Ew���0���5wq��P���j$'� ��e����\p�l�c�Y���F��y���V>5���|��k�}�I���Vuz��Ӓr�Q����ؿ�̠��p�C�\E���{�h�/���4��)�Tu�8�:`0�����V���ȑ�=�|�u���P���dݨgᖗ��Q �B�.¦,���:�[�,m�Cku�A�~1b������B�xvN����Tq%`i�x�WDX�'A���_~pJ�1�+���=��
�.�]Ѐ��{uP�s��QD��IY<�*g�p�Y7 '�zFI1VIg��k�jJhF}q��8�8����#ON�x�õ�
�"
(���f�v���~���V�f_��ʒzc{X������TW!N�ep�:�x�Oc�22b�5߳��/���g��lY�c�Ğ�Ĩ	����Ҍ=��۩�tZ<��Ir�+�HvRZ�Pʁ���d����$/��~�⦺���`��<��>4a���:�� G���'o|����ՁXv��/�"e��p��5�Gg�>�a]%\�љ�qxh�BG� ������	2T��T��P�N-���7�d;�EN^�|oOL6j,�L
D��ol��1����W|H���f�2䣝ʄ�:N�g����!�Q{//3�\�s�?/:�"���[`�3� ҉��HS2DW*��-c+
Ĕ߹p��I]���9���f�8�D�����7�&�K���0�'�;���Hr=%q@�h㾗O�G���T��W����k�K���Y�]azq��G�:���2$�@�y b��Il�Sh�b���!Gis�V-��F@ʜ喍(+�T�\��oa$\Fj�����_�=|PhA	��(4B��:!���	#��͸��C�KL^� ��=>�y�d�}+zm�&�_J%��C$��{|5i�b"�)*j:|��hCEB�������a����M�����2���r�'0�Y&�IYJ�r��㶗�q��{:�[kn�TO���>g?�{��'��$��d��;��ZS�j6�?WE�%��.�;B��qo�$�|���,Z�����ف�f�"6a���1m�ax.��d'ck�H:���4#}���2.0�vg ���$.AlZ�^��a�.�Lłq�F��ƛr�c"؆%�8���h	�k��a)}�!��E��V!�h�&{U����
��2A��x�C�J� `�b�=��a���TR��H.�яۋ[�O
[����	�Ju�g� ����F~$cbԾ���M]i�hV�Ѯү�[q��]�CA]U�{&n���q��M�
���>�O�C)뾌�<���kg�v��b�`���d8l�[�6>�i�ҏ�ZlT���]�����<��]�Q���Е2�Ր������c��>R9!����P��")l������#���jUc�
{�� �\�PF��%���I��ٜ�g�2� O�%y�8Du#��1�0�	av�O��%�%�o���H,�$���H��3��%�fb���u|�w'��Zr��b�q�4ot�Auٚ��D�24������2��څ*C9���7Vi�[��&	9���zכ\���.�����c�~�x �!~Pp�[�m:lӅ*.���L�X4���r�e�å�S��P>H�d+�R��G��w��sfG�n�����Dhj�h%�p-���|d�wVuC��L�Dt���%u�.}z.0<����˔��������
#�(۝������`5�u���.���I��c�0eIn؜ļ����))�E2��@(��]�þ�-��?(V�P�����t�$\�;�y � K~7�1Z�=+�3h�a.G	(������uG�3.|��DSUsE�������nkց�욢������!o�M.�v��PJ=-��	��V�N��@S-�Q�1\�r��'�A2q��L!x��Y)�g�y+q&��dM]3)���P�Fş�T�V`o�������H�y}nlw$4�����%��BȔj$3��m�#��^��NZk�{&V�f'�UjX�x��n7R��;�+(,�m����eB_˲��ۤ�l�{��4'	�#�R�t��S�+Z�-�]0����7�1����Z�I3_��P ��S���\ـ�7����~����V�ѥ"�=���XU�R���d^���T{��i���{�`����N��zy)�����?]�$�`�YU5�b"�^���k�� �nG`/Ī�%pB�[F9%Z�	��ւ�[&�)["� �ĕ2�j�̣���6���t�eH�˸Xz��_V��"^��Si��N��k�%�ѧ3S%��Q�*W|�ބr����2P��CO�Ά�X�m�O�L�E�1�ß5W��fq_�K}q��F?Qu�h��a=v.�J.R|�j#������,.zH�\�k!��y��RC�"p��,����[�C��؍��w�[F�9���`C�P�c����s�����Z���g8ڍ).G(N�r������� ğ��S=  m������j��g17w��C���=P.C[k���;!��-�X@�mZ5�ukw�$c�ܭHL�"�a�19�M�?��T�3
SMO��y]q���W�~ii����gp�@KB4�K�8��D��)����tP)��S�Qjwo�z% �6G�@���e����N��se�3�S�
 �I<vn�	+k���^��f���L�e�xr�҉��b|�&L�Z_�'�M����t�fUg��;�?�G�o��[\�H4)�<�|�Fi��̍V=+8�ر�m�8��8��\ ��O�2T��(���\MV�`6q�?��\,�h[������m�����x�D1�b3a=�^=�!���i{ִ�
���v�J�iC���!
����Τ�ɇl�?���U'ti.}lE� <�� �?5>��%y�h�v�Ő|i?I��$@B�bf]<�|r�gםd�0�
����r�d�ٷ2�G;ѹ����L�#+�!c�Nn��E�[����zS�!�I#�
>�4��s�.�m?@��݅�.#����-�O�6��&�f���C-������(�R�����:4��
����^�I{;<=|���ܰjm�;�E��H,�_S�Za�|u��E����h-��2{�~�m u����V���{��Ҩ���;WA\O?��Y�y�k��9����pa��x����]b�3nְ;읆�cl��Z���T�(<59X�Q3��E����H�%�+�m��coa,��^�v�&P�ZN�(w<��g�js��m}b0�����\/`���7��б-���W�%Y��n<�!m��}���x.���DM�ȼ�_n��DnO,��ó_���}Z%µD�!��l�&�U<¦rU�)t��@Mi���';U�/̵�x!~�������q�ʵ������ V���O4����Y"������0����JU�����G���\g���ƶOyl`���4�T�Q1�BU(��atD�t�TW��1�P����#"?r >�վ��MZ�Y��qv'��"��J]6ǎ:B�΀HX|����)��kt��ߨgF��@	o��ĝa��Q�^�L��>G��0F��+��_`�� ���~<���%%�j�c&�v{�F��5���3�ז2eZ��ӗ\e* ��>
S�b���cC�Q�=��J�Ϩ�Ƕ���<�<��hV1e_�|��q���6���Ϗ�<�ǚ�'o���@���6��qk3�b��V3��gXB'\Ǘ$"������8���M��S���f�^�,���x��
�yK�\�o[j�.���<�)����u<�cN�vI�p���٘���>�#F $e�3G��N[2�܉�-:1�y]�H-�$NQ����I6ElZV-���)���E[l{���3��������W�����:�h5ǰ~iƵP�.��I�X���,EC�ꭷD��.X��1�>�т-�߉Q���(r��%$J��K׵�ٓC(4������}��\'�Q���C�YJ�M�C+��
ƈki-�D�ڸD�U�
~L}%,
>5`\�{f}�����&���t�p����k(+ S�s��Jb�ϐ|��
�7#c(W�1�/Y�+�����Y��#�E;���>`f��s����E!
�V~����ș�Uܭy��=`s���F;�M�0���aq��A�͆	:�ٕѿ��o��� �v(��[4r�:?�ͅ�y���wd����XD�~E�d���iR�ͅ�OOq�y���X_""W%�*/ ��O���C�m-��/�biHhg����k�+u|�,-�)����
�Y�ߥq�t�]���J�&Gk��P�I��0Y�,h0��ϋ|�F" ^Q)Tz=(�>���|�C���6O�@��c��*�*)3�@{�IN��xwZ��y#��Щ`���xBVL�I�;mKG�kmc�� &%����?AG���[?ݣ��+:C���煫#J��HP+�{����N����
ke�.�ʊ�oÝ4��몐�Fݱ�9�jD2�Yv��xc��w�[k���Y������[�7.�����ؤ^�E��B��hOU0ڞb��Mu�t���XKCdF�n^�˥J�d��h~�W�N`�㥯s��R�L��!��`r�m���9���<�B49��}��%��z<s����O.5�NU[�ż�pĈE��tcE!4���R�cs�U��߄}{������U�L�V���T-�W7ч�8��M���6L6 �hl���PZ���Wc�O�+�mv�v��k5��&U3ͻ�3aI!!0�evN^�+�f�;|�� �+PIĔ���z�*�3�~x��5����名_��|����� gF6��_Ep+RM`}� �(6߮�.Ա��yB��*�"ju�VK����:ϴY�U\~�ӛ��Ț���m
�?;�xr��P�{�yH�b�G5#���#���C��#78�܆�1b�: �x�~=S�A3�5b����8����P�ufA-ւ_��^���1�� �>g���q�4%X�8o��?�O�O�ZQ"n[��^;��yř��^f!#��7��k�E9�n�:����Bd`���[>���Ǒ�vL\�=ϊG�鉄�]�r��Ivu�:����׺�tH�n�М �S%�h���C��<�ס�& sǂ	ɳ]�(�L-��B�"�S2l'ؔ}�!x���_Z�o�U3�gDG3�Y2�C6���\� Ce�faT�Ni�P��\f��	���������3݈%g������*����L�8�#:��AY�
���8��1�]�IP���M�]a�������$�o+��M�Wqvsfݵ���� ���,��kB2o�}�u�B�,����}����^n
}���f�v'�r3�2��H���~.�g�6A��:�,�����J������a\Q�
w�G�;�!
 .�y�&QU{�&�t	x�)�4��03����@���8R%1#��q%���R�����j�J ����=	���}�mi��*D�"�������k�� �fEڵ��4����r���\��u��S]�pq����y~�U훫� ��-�Û9�ALE0�q>���������5O�'�69G몾貺�Tjh,:e��"���/)e��iV'��t���I&x��W���l''C��_U��k9��q���J��Aj��һd�BD�!����� T�,q��㳓b%&��7�늝4��ns5�n6��b�"-ϒ�,JYo!8\�����N'���3���
R��;�,��]o�]�cH��nw���E���%��xy�����2����D+4���QT{Â/��"H��ۅI���:���4e:��7>�uq���g��ڃ$�c�p-t�����*=2-�LO*�,Q�`l��b�J��;LM�	��h֎�Y5�� �xL���-J,�*�x�n�.~$�Cvl@Q~怙�Y�P����A�g�<�5ꉣPuzBN�<�3�!-����@�^*D�x]rܐ(X����4�=#���� Y�p@�}�On�.qW���>z����@4S���aF'@��q���^����ç&(�D?�U;Z�Hw�<���M��g_(�1����N@��j[�Ȋ����A��؆A|"�s���fsRD`�q�������r��*Ps���g؅�hV݊�����W�������C��O�dNhI|��W��M"�:�R]Vqn�G�%,���h���wi�.��!�i�ܢ�Z/d���3^�B�h����Q%�B�Z��'!]X�H�kx�m[�S拓嶎��F��{.���؉��#�"���T�.��E=x��Z|�>;;}V�l��;@�� xB��C�A�m�]�{K��A��_H�P�ͪ���^�z�A�ʞ����D����@����ľ�xZ �,����G7��ɞ�.�%�j�*^�{v�>��������.v%�#���|ߩ2�Q�YeW:��F�779�C�'!�ŠH���q�!\��"�T���E ,d�v��͆p��K��q�����2���r͵����G�zv�q@�M�+�Ei��!tM��7˘�{��<���^͕�س�f���S��0�CV)Wˊ�>m��[�fe�@ul��7<�N��\�bdQ~p�Ľ'�c7z��}/:NKm� QU�wd��9��Y���9YJ$��<���4��&�^RP�迚lҀ�!��p�⭽�h�c��`
�?��L�6Yv��%�p�sL?��ќ�fbL�c�P�rL��N��\]v�p�ؕ��^��<tc�(�+����h58$��#�PW�c�ku�D�w����њs�h���'8�p9���x���d���������6�e�턳:
ҫ��l��[l
z�H�`+�CkU�����|�KK�18���&��k���l���/M���!g���2����.�Y�!0��Gj2��{0��:DTҬ��O|j]�rOj���w���w�f���f@�!0ri��!D��Vp�ڋ���h-u��L�9n0�&<�Cs����jM�yG��>�6�w)9���/�S����}��AG�b[K�OFB1��yFS�R�
���� ��{�eܟ�2RW�tG���࣠x���?�<��.a�gWZ�L�'%���Q��q��\�KT�jG?5pD1:ܺ�?��AE�-�)��W��*a-�����m�
��:lD�pw8��W�4�(���׋�Cc�W�^���6c���Z�@7��ұ	mc��Ƀw�'/~f� $�.��˻����;�]�LbJh�#C�iFF~����"��Y�Ϻ��N�(~�L�"+ꦶ�rN���=W-?s�d˘f*. y�H�^4Jً��������}��ye]�	#��nl]�F�=&�&�Q� 螎�x
2�+X�$��X�����Ww�FY����}[-�|�__8Od�,?ƊM�7��Ǯ�mU���1��.��E�/���˒�� A�|�'x!��i6I��d��z�&=fAA>Uʛ�(�	�����za�.�<��c�ȳ�᰿�D�B-�E$����
�-8�i2�����R�l� ~5g�֜k	Jq��<��j�RF������Wҕ�n�_���_lw-����q�Q%��ŊP?�
5A��II֓H���mY[!�ZI�U�S��y��2�>��W�O�ۅm�
[V(�jeES�����a\�.u�R�]����J
��&�s�-a�}�[U��1H�
��/����l[>Ī�k�K&JF�v�lX�N8w�l��=��gF��$y4/�*i����b��p��}��y���
y_h��u� �Vf���l\�m~�B�+�
�������bW����
�Ƅ��YZ�uR~P��b;m���ɨX��#װ��K
�˖J��d���'AJ��'���`*�u�i�\Pe�`Q��I �����*�,��}t�5 E#,�)��<�aI���4�M��gT�����J՚��?��50�[ó�>�OWl�ФV@�p?fg�t1
�&�唒}������C�H�0�.��mM�x� a���93F^��Z��sQ)h�-���B؄}	PM�d�I���mOe�W����fXV�˅���Ϥ�L���X��tQu����sL�ǥ7����[�2�#ӄ�j��4("��!�|\�G�� Q�ڼo��e�%�^:y���G�s�Šڄ�#���#�O�.�/�N.�R��T��A/.'Yr��Į��l�טj�Lzj
<�5���s�3I�_^Z�)�ӽ��=�L�FNL��C��J�o3%��Jee��U<^!
�n�%ξRiO���gJ�����A�X{���y�AX��=���w�w���!�WF �4�maY'�[��h�+�U�r,E����u)��C-3�t���c�kU�e�B�/���b(g���	��s5]JƱ��f�L�I�nU��	��}��ϥ���	���I���U�^;z������=@t�R�on�V��o��(�1��lw'��?iS筅{�{��A]�t�Ҏ�p�ON~S��������`�Q`��;c��ir΂�_���`ǟ�����S>�����(z;� ��6�ae+���v����[�{��9�����K�����Ԋ��L�2�s�����<FQ����3Xb}� �3z�o��|���aQ尢���q����TwK~��>�<8��n�<�W� �8U/���[��H�䫻W�U�H��=�i=K���7�'/Lb�)���(A'T��t�J_<L!����uq�����U��D�cF���'�����Ja�V�C���L#�y�
�b>,O��v�mp�N�	P}�{m�`&���
�����S��ыsç^M9�EwO�1[~�W������K�A+���6����:�-�;��OE:���AA���)�CԺ*�?�	aH+,�p`x��.��TcX����G����,��F"�ҳVFq��A�U�O�����3�崁���T�78���2!W�xP�O���ύ,;����X�S~�
8RC}j�ȁ�����a�C��h����3��G�E��Ӵ��I�7�6�[�ξ�ٟ��S�k��DO`�����u�U�&�@
���Ԥ��� �:��/��a��c�#T菣�.���xz���}gHOF�R�-3�Jl���^������Sk�>�h��`1��ןMN%S���9��?����ցP�T{�a�ߗ�TA�n��@���1���(�_*��)�J+g+������U95�{�^Q^����g��]�7�*iQ��_{�%6d͙�>)^�HT2��9�\m���/)x�~�l��LsE��VᝤYv�^����3K��e$�uVÞ>��ozv�!���R��88m��3�Ȑ:x��͛`-���ѿ�h8e��"������eo��|�a=����u�����e�h�m�:�*�3��K+���@��0U��O+@EJ�����]7;W�z�PZc���c���ʼ-�m2�E����fj$��[�s��PF�q�h�RJ$�@{Mx�7G6��8��qDM�^���Q��I�D��m)<�����Ff�כQ��O�-�E��nO	�e���2�1�O�zn�&K��<3ϛ���Ov�~� �z/K~���C9AA�=���j�q���-�Qoy�H����3P5��ǽ���\���7�_+��[�����7�CO ��G����)́x�4+�W�'��j�-;����<�7��{j�{7���dl�����L��[��_
��%��-La�ս9�9+D����m�B,��3L�.l�<��R�ݭdh"�7�V{���,w���NÜ��v\�������D�; �F�b�}*��(�I���I�)k�c�]�3�������9�����O��h/���O�R���Lw
D�3eo�G�
�-�3��G����~l�,�Y4�3�y�������+ �����?b���b���.qVi~m���!���M��@����;h
�S����S�p��<�r����?�2�6�D68��h�vg��ʳ�p�6<!e8�Xڕ�@k�0�3x��mu>�f�X��Ga���,ɟ��B,*ͽ��(E���/�Й�6����T��b(�$�!ϧH!H'�d�]��;I�ɠJw1���.b���Y���3��ޮ�o��]Nv ��w�vC!�s:����E�!S6�mhvjX��@���@ +%2MRȽ�~����~�#�k�J	�s��H����~Ж~�(C�v�ƺ��<����a�ګ[���:�r4�w}�G?eG%T��P��>x�+ݑ�䅡��b�6>���ۓ��.�aZϞӲ܈�Qn�^�W4&�K9�4}]�ĢU9P"��XL���]G��F%��<l���C�|5���c�E�d���At��{9�tP��)|�9������֪��	�!��t�d����zyF\�g���,pMh��0A��ڧ�`5������&�g&pD���>�0$�;X��f$Y�MW8=�>����|�305oNi�ߟ���n�UD�����e>:��4�Sq:]�,6�t��֗oDz�Sf;<�rhھ��0`ILp�!��֗�r��}�G�0a��e��,`ƸV�bӜ�q*�{�ϼ-~��j� V*K�U 
��f�9]j�7�M��'a7��p+jr��@�H%��{�3\��"�Ȗ�+�Q�z�����?a�Kct���Ƹ}y��2�t }��nAc��3�G�O���]�y��KQ��l�� ��r���a_u���@����>SdU'(]ံ�j�Ӡfl�0�f�覈��wUc�q��ǆ0�h���`͸@��ߧ7ƽBJ����\ ׫���> z��}����0?���6DKL�v� �.��;���8�ѳ�X2�k Z��E���z��sM0ks%(��_8O�8@-\6]��u�y��+l!e��ĵ�)�F�G���(��٧>�����7���bT�����
�^��0\����[T��}�!e�/]�d�]�L�.�y��p�5�/�䎒�m�L0����聒88@�Đ >��/�z�*�p'�����H*M������%�჈aR�Nms��i�Ԫ6�c��w��1�E�sv֯�^Ǔ�,�1�	P�S�a�g�v��
v�n�]�n�y�?�䠿a��(��̜=z�A�p�Ln�קWʐ��}�%�yw�Dr��p��9���%e(�����{+�M�L�rl2�8�WZ,g�8��<{�9u?m��Q`c
�Y+{H��}O-Y���ƒ���v����Ϧ�A�_t����,vg�-�@2��n&�[�Ϛ�G����*(9�iº鈎�t�!/:�$�eϸ���'Mg�q������^�����%ĳ"��402?x)�[�����@��U��Ϫ�X��B*�2H���07���j �cna �Y�㕼K�M�e���ڣ	}���G��=��Q�'EEXt݃Ҿ�
������6��IZ���,b��Ŗ�B�[.��[�2 ���(���f��X!��qHɰ7d1��Y^����3!	���U|�{y�8�3�gRuh�>�e�t�»:��iJ�ٻ,��\#CVns0*�wg����TFơ6�)L�^8��))��$��?�|�f�)�C�T�A�0�gd�����1G,��k��w��2��Jӓ�����8�
>�������VD)���F�Ctd�����ܵ�7{ΦH8�k�q�l>!ÞQ�Ⱥ�l�B2!��۱�!��51�S bn�DPe���֚j눒$���35������p�h� O8v�~�+�ί9�Y����V�f��~�N���J�q��Pϭ����x���c�cR��$�&�\->��C��r��!g��ք�au�i�uX߬�0���u��ˮ�������#y�+��q���*��/�g��?A�UX��RG�A|�n��
��\P��ޘ�8��>�6)�	r��a B�0�+���Ct��*e�(\�W�iJ��:��p���j�Đ��_��������`��"�C;��
"�a�tE��*/�������G���V��T�Rb���o����ච�/(3+��~	Ҷ�η��(9S��.�Ʋ�z΢:@)ꋲ�%�f�����Rއ�I��c����nT�sN��Ӑ����l���O�Z��8�
���5�H2�L��� ��ZjO���O�x��A���a1��c#�@e�ӵ���˧��=��L�4QE�����}���3!�3#6sPc[zA/v͉ U�#6��
� /�����d�H5�����{�i'v�ϗBZ6���o~k�d�N�5[�������A ��a;F��$�'����]ꪁ�\�Ij�����,ֳd>�5��oQU�K���7���&u#�\`$��R�v�}��=3)��"�q;*�> �9P����5@�-Ld(?����d���/�.��T�2KPt��>�m�pY���`3���d���!�)��� yk�jG�Y#�s��+�H;PO��燮hl�r��Q���/�Tw��A�Ѭ"i-!l�)���B)/c���������00�
�J�E�Z�Q$W���a�Zv���ëG�v�
�`3V�B��S��QN�� �щ:B��J�ț�{�:2Ț�p3ȣ�+�����{�S�v��+�`��S�,�
��5auʊH��j�����"��=�,sNk�b'�F�ws;p�ʏ+9�}���I�cB
��<p��)A5*x���:%2�5�*�ᚏo1����O�����Ap��6�~tܓ��覌��,11	+/W%.��p~ �8Ez齉��i!�t5�1�q��w�y-���a����[*{3K�H"7���� �P���1a�����?}�-�9���P`�b�'�(禛�m�\8:�f��1��o3*�cO��k{�Ar�_��V}���$YCXg�Oу���	��dMw��u%BR_
�sz�RXn����������*h�֫�	87�W�E�ؘ�.��e3E�Ř��R���4��8]J�9.]�b��F^�Z���F&4�+i<˿-r�b6��D�� #���H����ϻ��?2H��@���JG��Sl�.�����iq�6�Q;�
�,���C�����׎<�2%��@�$�$G�)RC�q�����4���"k� �ueE���EAn`F�W��M�9\W��{L���2�1u���
�#t�&�0��y)������,������Ƣ���� ���z�d:��a+dxe��Z�,�H|�rHj%�+��w��6���@H��n����(��A;�ϯ�K��-M�{�s���X��'CT"��/��$4���>��	���x$$j���ӯ�(垺�5TI}��w�g���GƼ���@"<V?��������'ͰX�T�}��fP�^��FG�H�d�S�`�ZG�|������%���X���L�?�A���VVJ`�u�P�����������_��T�w/�'~�Y:�c|UY���cP�w�Ƞ�ϒ\x�A�[�$z�xz���i$����{ШT���U����wu&��K�]rQ��95/�r�v2|癇�c�L�j��8rZD�&U'��auQ�G��c�I�2ՄP��5�-,���_��v4�v_�{}�d{�<����}�W���)��:kIZfM���Y�$$xl�Y������@�uW+.�PtY�m-������])�3��-�l�'�p'X�2A��"���~(�|�3>�<	�#V��Yܵ|w�ڻß��*�%��o��m�%]v��7f�,��+p�%�=Y�W���r�Lz�d��I����-Bd��B��B�Y���(	�ql�6zj��6H��^ؖ�zĂK4;�V����D�B��;�'��b�xE-K���y��`]8��6��z���K�i���������n[��f2���8�/�1fV�����9W]C��>Šzt+��l�co>��i�?�l>���Մ>��㬳���'=�{*O�ky��������TJ�E{��m��m�<�5��~�M�[�j�1'7��MM��q����-�.ч�o�(�xLPe�a�|kB~���К/���b@������eЧW������;��[8S�J6Q�7?Z��lZ8�����(4Fy�C6���pkbD^��"�w����q[�"��#�t�t,=lj�	`%.���S�6@UH��Ɋa���1�����+�zW�Q�N���͉T���ޔ��	ea�xy��p]]������ŜHh
O�����K�.��a�P�ދg)P!���O� ���b<oRC�g��K�&�h"#h�o�KE�2ȅŬ��)�e�}7���4��n�ҝ.��,��wg�ʰ�I���}Y6ϳ��3W`	Y�,�Z5��Q�@yb���h�����B��]ܷ�@$;�
����0��\!�'?B� �4��]pa�.k��2O�|}����P~fk�p:w�Av�D��y	�n����4�߀�t<LP����_43j��;�}�z��z��7A f	���J?5O������f&v<&�E}��r@�����?�EZP�gv��Bal�O���A�2l4��SG�:4�1w����{fb�~ٔ#	V+���mK�l�>.[�*gЌց�@��}�|0�:D�,�_>�hp-�,K�	MdÜ�C�xh�/(�����(�?�$W�A��j���ƽȯ6�?��	��S��1r�����I+Oh���g*�ҷ�㓵8�f�(����O�C�S���hb�ݑ,�T�i�w�V�l^=90�!K�Sd��o\H�8F^ݙ�>�+e�M��vo��Թ�[�RCvu��|�c6d�V�&�d7Sd�	��ѩw�+Ym�����0ȲT�� ��upyW}n�R�u�J�N:d��yH���ߡiڃ��8<�-����ZЭ�n��],��hK�y�p#SE�ם�Q��,�6��S�����	�	����5�L�CI��}|)'|N.T��#M�#�w�G����aZT˺�.2�`g�H7C�W��*Ն�n>��+���u��"ΏJ�q9!v���B֔����ow�.�E}�]]��A�q%�o̟3w X�B��䅒o�4kۤ-�_�#��ݶ�L-	�%{��۝p��,QW�1�3�nG�X�(���m\�u��	N p�s~[%�N
w���P��Ğ�c}��}���G�9�����jx~r���N���
j.�eX����܇]Ç��0�y��6J>H��iZ��N�=Ѭ!�LI�����$�k��N�~��s�y� �ٌd��+�7.�oXZ�G[��ɇ�T[���$o�v5V˜4�~$OL!Bi)��3x���e�ig��d�U�l��t�qQ�O,�����/��6z�}��-h�b5�&\��0�kL:��
�ƊyEgg"���U$�1Q�����q��@`�l�[7!8.nL^rK��6>���D�!�����(m>c�R�����S��ʥJJc�� �I<`j�ꓘ!��pv,�ӋI�Z��fi��S�!`�u��L�@���lddU�f`r78cS�S��R\_W_y���HqS��pJ�9m+.L�x�`JF�*����%Y7A�@�U}$3dl�V�[���Ή�.�!����E	I����6����: �NM��|\���h��s�7|�wcK��Oã��h tIų1��E7�eP�Ia׫�k5���ɯe���%�
���J)��7Q
P 0�o��6�A�z���i@�`�<���A~A���tR�cťGƛ�:=&�O�&�(�hd��o�Ӑ�*�l,�x���R���4?b�!�JVC�†i1���g���?,u�˅ �~#�S�*�/C�]Z�o4$���޺b���~�t�{T��__�/doyG�ԥ�λ��9����g�+�=M7�e��h#�s�c���+��:2Z1R��
�C?�1���O%CP�5���F�xX��De�@�ܮx�ԙ��D�2y����fE�>��ļ��E�Gu�ۉ%	z x���I�f�3p#���%��{��,�7��]?Yn����Q�RSd�5
{F�+���#/��/�1ZWu�4����+�"!��^��pm�1yO��M�O 6��X��0��zR���S��xG�߼��4�N򈕪8�(�&�gꜰ]*ݫ.��F���E�X4��:0t�ټ	&�fn0�1�%@GUP����^�%��9 7��O����]Ay�h��_�9�� '��z$��^r:��X%��4��X���y�̗`�S����U~`;R��l� 몞k��f,����L���,'� �sF�VJ��hy���|��y��� �&<�t'9�	X�$�R֔+D���i��n��Wߜ����D|��WM��U�ܟ�`����rc���zU���`��p�	=ׯڢ!�m����Np4���A�NB`u�����-/W�f�ؗ���t�)~(�}�Y�P̤k&mw�z��4�+���Q0#��&R�J������=Ǒ= u	����AP��]���(�p_. ����kE/����b����kSېK���]emӱ*`ܖ�p4���C/H#fF�M^���X�^-����6S)lF0�њB�?�`i`��0�D�PHws�����.�q����UR6�x)��t�:,��佫�� ��,�������I�r�n��3I
+;Vl֎�GS�{�@��K ����gyA$�liF��K�-�mo���\��r=����床Q|�|>Vľ�����ɢ��v{풚�[�;w#���h�{�\�
�����[���d�>Aߠ�/��\��U䜍u�eǭ��TG^��r�a��j�K�h�Dۢ�bz	a�����˒ �G�W���d���3����9R�\�eS�-�|��pS^4���B�t�&��l[E����� W ��
y1��#]���Pgl�k0=jc%��	+�,Ģ`#Ϛ���-EC7�K�s��:��"a��t�y�
�Gǖ�-D������������sʈ�.�����Zv�5<~�y哪�ր�&֐)T�vPNc��vL�\� ޛW<�����5X�B<As�hp۔8��%-QpF�E�"b'Jc�'�8����X�	 �Af���T��d^�a�%8G��#X8���Z����
Z�A��W�mS�e߸C^q�i@=q=pw�C����-��O�i�$�K�Jۈ�!�����!��^�Ck���J���x�P"�o��?S2���d��
����@jS���T�i*�l�.Gd��Nyi��'Q���׍��3�'�P�1��fq��	�0�����|L�]�(��,�u#X:ut���''���� a`��9�7<�r�0̹����q�x���������eҀ�J��l��5!�+�R�m��W��i�� ��IF�u�+�P������س���o?McLz5t,�؂�Փ�K�ʕ���j�	�j�=f &o�֨��� ����m���͐�
U��R0�c!Kv�J� 1��tE��Ӳ*��:P�T����� �:īS� �%�y�:���S�BN��yq1�N �r�P�G	��y��/�]=p�a:�����������h�N@^p ����+h�"�ڋN�d�dZAp��/(�)(�����KD:�������YX�7,���͏�
�i��Z�<d~#Hy�]�9�\#w�T��$��L�\�O�!t�?��F~��*x��t�N��,XC��2_�}����0ƨ�-�i&�\N#5���犗��W��F7�G��|�cq[<�:F����P�@$rݪա��!t�m}淡����2X&��5�˫c�\�d������?s��X*��`Ar�*`����(���;����j��
�Ø`QI��w 
���(�,�("G�o���-���08B���.X��*jP>�7T����'���~�V��+��`!� �*���)���i���)o�V@��)�0Ò�S�Y��$��yL�	l�Wp�:A�@�R(��#�:f�,��SpЂ��Iz?�x���!#�q�C��RXf	"zh�9��GՋNf�4�۾��:��2�Mh�rEЧt�>p�D����Ŏ�_lbU�4Q50@]3�c��f��=Ke����L7�.�l�������qut�xU����dOfUgf�(�����!J�A��\�oO�>Ś�j�i89ZD2��:]H���< �A�"Y /��O;�#X�tY��Ě�G	¿�o(�Z��-�0؟.Q ����eaY�lƺ�����<b�vUo;W����5{��/BEs&�)%���s��a��q�~؊A�VbM'����Q����7v�$����ƽ�:�3�~��R�£�JW���;)�6I�VD�Vn,n��3S}v��Ŵsnm�q�`�O��xأ�iRX��Z�^d�&��KpY����`y"���������z�-��-�E��zUFC���`ҽ��0�;���qx��%�R}8�a�wx��
��e�B�L�s��(�i*՘��5�b-g�vq!p�2D����}��;�&ڗͳ�.t�&�'�R�$������H ���9����m=��-N��w xˤpftڪ-^ESj��|:�V%��g�o���KA��ua���V$y�*����y!p>��?MD�%�����]@��íe���v����(�,�s��O8����p�-'x[�m�4���Y���������`&�f�byXT-���z�@�U5!�L$�9��*���_��
�D��^������:�΁H�	9�l�� ��@�Ĕm��o��6Y�Q_����=Av���^:����<",���1��`i
\��\6�G�=_��,�ê��I;tm5��X.�b����{s�����Rq��N��\U������q����o�*@Y���:�qÝÄ���G?���g�ƅ�/�Kg�\���A����
 ��h�I�d�jZ�
��*�h�QO��g������]�.	�dbRݗA%4&�˺X���p�iO�u�G�&�m��@���g�?���}-{xfm���؏yAk��?o�;����0l������oۥd�nf�lUw��K7��K܀��,?=ڹ��I���<���s=�;���,��?��ʫw�V��S�,��rI��� \7�D�E2����|n��V��^^���׋RG%Q}%�P�ĺ{�q��]����i�w>y�J���+Z	Z��l\��[\��E�(vNj��H�O��Q�"E���Ĕ�]�rU'�eseB����/~|��(ۻ/�ژ㈲�@K" \%�p����1�XI
��T  ���R#�Zgr��lR�s��Q �Ak4FJ"9�Gr�Rwf��U��v6}�f��@V��T].�u�}�ح�4M��v�:aZ��/+�P�&g��U�n���m\�v�1"-:R	����;8��;q,R�����������7��BF4mD��p�u/w���X�.0�V�V�8{Q~�����-J�g��LnxH��� ��,=�S`�ǒN�a�i]U�B��X1p�K��#�>�S�8_�ݨk��~m6������>܄��a.2e��-��ED�0�ί��.V7aE�3Ъ��[�kg�R3Z�dv�vr��؄k<�1��s���P�s���۶	�H���=3�D����wu�T�
}�I�������y](׵Z�	� .|0�mx5��r�_@jX�͏Y+HZ\-���ŁSS.n�i�	�`���y?�Im�K
�ָ���`��]�Iu �ӫĦJ��!J4��FZᳪa|�2��K������n�C�L<7�S�D�W��P1�|�5/C\0�*��`P~8>�!�����*f�`r�l!YB�/h?Y�}� eD�VDe�߳�%O�C�s�E�+a=lB����"	߸W�5��fe��,���Iy��A���v_���]g��9+D�Pg)'�X��ᓅ�l��t,i����	�@�R
S=�ᦝQ��)t)��X {�� ��yw�M�P%/�u(�ީr���ˎ��3�.U��I����������ôB�7�B
�Pu�u��z#�k��?��IZn�b�+I����(?MW/*O}�"�-�'v'��	�2��<�Lpv
��8h�����A�F4��>�YO��.���MФ�Oy�E�����Ec	}�*��	�]G(D�E��[�A��(`�n]tp�辢}yͲޭ��+e�|��Lcɒ��QF?���=�,�T���pcn�ˢ���fu�f�$x��oy:0ѥ��U����^!�_��q��A�Z�@b�{2M�i�%�b��2�����V�@-�)Y�}����6�~I���p�;̗E�%��m4���b�Δ�\��J�܀�������;G�����SC�S%���i]��20z1@��D�����VdҐ�����.M�^A���l� s�@��X��2��f�@��e]�6��Z��@�n'
�XeBZ������߮��w��� }�\��2q|��%�
�@�.v����]{Mޓ;Ѧ��i�H�~�h�ߙ+ݘB=2wXiVȶx��?��+k�Ep/��Ty7Ä��=��(����Lv�~�T���zبy;g�(�F�A�����{C�=[����m~E;��Z-��RKg�w��e4z�*d���y���+ؘΚpw��- oU[����|�#��Y/��z	��h`���%F8<c�,Y��Ĉ��ضܕ^��8ܥ��I���	&_�[�xX�8D�6�4�XY���&����Q.n�0�Az݂w��WU1`�Y�2?���� ���|�-93)��:�䏷�?�@�$d��\?-��VÒ߾�hQq�&�7�IVoO�K�L�̰EfI`�k⌗�c�6�܀-	�w,�%�@z$�7
R|:�0�Y/[�o���Ȯ[�ɮ�E��>�0�f�����ʻ�"�OS�)/�5
�uK����Q8WBVڻ^���Bx�ޭ7�D�O.B����/���U���#�m�'ºE<�����ۼ6��Ϙ��Ő��@[����M;�yn�
F�)*U�v9#�����2FI� �G!z�f�L��-
��5Sk�//�ֵ�c��ٵ7#�v�C�F�i�x�B�_��Vٵ�1S��3x�!*���y!��(a���Rk�-�]=�� �7�".Xݾu*��r�M!	�$�/ބ/����!�C�g	�0�G�|�殆9#  Hs��E-r�sL�$�9J�\sdJ���U��`���	h4>����:��΄��R��#�������ƈ�Lw,Ip�h����4�GB#��L�����5�I����CByC��
'��a �<�Q�{��z|�Qv��aAI��ly��o���c{adQ���d��g�y�6�*R�hf):C��;�4X:p�w��%�=��~P~�Eݐ8��MVCw�r��c�k��	��I����?��t]���~G`dqg���Ɓ���@�Փe��9�$@���x��Q�`�oH)!N �g��rzIz���W�Y�U�_j��<�o��7�C���@i��\A_9Ȇ���Cd�`�y��<�Fe�B�$4΍�km�(��*f�;N��b^���ϼ�: �����f_5>l#��+�~w���TB��(յ�Ǚs�#�@F����~3����_rc��Z�H`��f�J��C({�q, )��l���.w'2��K��R�l���Kv�?��m�O�lHhI�&����9�0$�	6�p�J�N���p,�j���b�M4x������}YÝ��l\���6ظ�Y��[�(��f�I��*��eWY�}*�mN���:��ހQ�2��|�ɒ�R�{ơ7$�T�$B�J���lE��O9�E�n���*M8�I/V��6E"��R�5m+�/F����b�>Ew& �"�2A����(�-8�~<�%��f�5��L�l�AG�@OP���G׺�	�މ����E���n<�}���)	�0���'tm��$�*b���C��d�(A8�?NE{��ˠz��z^��^�(�ؑ���e+R���v�}@�o� �2&aF#�W������>T��I�_5*�>r��,�9SG(R[t��Xn���. C�3?�q���F� ���2,�"�7�~��/�F9�sdK��dE����a�b٫y$]�M ��X9yCԦ���V�7�|bj]���Ύ��jC�=�gn:_�'; ��g�#$W�@��Z�U��N8���0�K`�GI9�X޻W�Dβa�ǐ�պ���L�� >-y��`�S��{���P�f���RXz�䥧�W4��X����Fi�񐼾.i���3=I!�}Ƀ�[mW��tI�޿���L�j%��ȃR�4Fz��V�Zt\�k�
!��aƄ�~0/,�Q�j�?�����f��ɉ�c��bv�[-[2���9��'~���\��O��A��P��J�*�=���g"Y]r��v����Y�_��a\O1��&��A�=K�=�A�gDy#��AR�}C��-�gJ�x���0����O�qK��輰���DL
��4���[�����L�p� �8_���j#��=��W�����e���4�fS��:�[�|eX��7o?���6���[�J�Hzjkﷷ�}=#+n,G��<R�0M5��T��g����y�A��xY�>�r�+pI|���+BHE쨠���}�A�̠��X��o�~�;��� M����hv����9̄��4����>�V��C���C�����L�5s9Lں���_��W`OMpశL���;`O��4�bk$_�	�U��+{m��Q�'P���3�F¾���;Ze��р��G�H���������I���j^��ٯ*d땏�U��Fc�&5���H�l��y a�q��ȃ�ڶ�"�Y�-DG�c�t�H���b@��O|�T��)Y�~���`F�(�WN%:���*�e����%���Ȅ8ǼY�~�>��0�w�;i���*@����M��&��;�9LUo%v�??�ǵ(����W������ ��	�W�o�����o��� q�u�t�C*���=\�d��G��^X��68{�\ �e�N{��^�Ϧ�	�"�i	[(�5���oʴ�.��J�+�˯��/��zL�ڮ|��`J�B���"��V���M����a��4g<cQ��J�O��PÌ-ZF��8�e�l4�$˅����_JBֆ� Ɖ�,n��xuiҘC�|�M�ܼ@>&����B4�l�����= m�wQ���HNT����r��V���E���(������2�
��+�|�7"a�I ��6V=��q�lVO?�!�s-r���L.'�)�Me�h���V���(,m<I�9�֜��`"�ĵN�+�S��
1�H4a˅�`�@���Z!�C�2a��Pbn�a�9�5�p���0�Z%����wS	�;t� ��eDY*=�Ie��.I�-��Ѐ3��3}��"|�Jw������*���&����0ԤR+��$�G������ZbS:e�#�W'�#j }�tMH��t��Q&���S�gSJ��յO.�Hd��2��^��z0���L�i�՗$��"�?��J��D:�B�nR���*�H�T=�xLc�(���� ��WܙO�(}�"|����[�ɪ��p!���r���&
w�uK����Kq�\��7�� �
p �|���+fV�R�oQ�����f���nh��T��Pغ.@+��_#��Z�/�r�*��R��}N�;)6�� =�B��;��(��D�U�w	�o��o�.�a�/f���\�z�݁��\7ɵ��iX|�%a	���z��xT�L��*�ɪ7i n��@=���t
N�> ,��ԔXɐ��@��U�*�����-�$tS�N���*z���zvB�<�s񜚶OT�#Θ�<�|?D�#���B6�:ī��7�.�/��m^ƌ���P��.��P�&i���v���}�������P�H�HL�A��]q�D.�����U!y��@�x�C.:�SEhE$B%���<R�s��j�L�1�\*��L�r9�l})~�4��ә�Q�l��ܘ%��
"��[�J��"�X{���ww�H���� Ȯ!2֝/�OB���D/�ҍ�`��M�O���J�������Zu��v��y]:b�z:NT�/U0���ն����ݼLG�Й��!j���8���]dD��p+�]MxS��%��k~�e����0���m%T��/�F1D�3������\)i�J�h3�y"��!�Bd�����L�DIOh��������O�����?�}�T����Qh��OU��a`j����Zӂ�?	N�����O�WDmj��4*{���g�R�n�#� �`Gx�n,�����DlƟ��3$K�~4��%��ﯨ)[����ۙPBQPٯH;#50Y^2٧D(�!�m1�Ct!��~�.���f<��oޓؽ�H{K���>�6�Jz:����w���.y�!�����	N�6��Lg������gu[�}�k���+n	*������k�ZU�	�8/)K��4�=����M�w��[���^��B�m���]�,��8�%R:��Ŗm ���"/<a�k���1�v����`�o�� ���${n�T�Td���T{���d+G�k�n�I�������6䢩��d����w9<s�X�T*��X���eٰv9�G詪f<%[%8����n���G=�l�� @�|j<�m��IZH����J�$;�P�Z�X|��jY�Ŏ!}�X�<���Z+����
&_o<-3�2�q�8��3Ԥ�l�ѕ��y/��w H�J���B�����"��[�E�SR6n�ܾ]N�4WæO9��M��ͣ���|@?���\�AW�Q������?.<��`�V�,c�u��~�>���'ɹ�^�/ J��M�ȁҴ���g��.����|��&���7����I��t}���6����NIo�f{[�wz���h����-9�Pv�����8[o[#�,z����2���`9�<瞇@J��͙���U�jVϴ,D�NYж�#�|/��^0�he�s���v�5o���EdI���w��v��+�q��N0��B��`>!�a������ ��v��C�}Y��(� ̣C:/��&��0QJn��mG�+���L�(i����znyV�]��>^K)��b�L�	x���Ut{�,�7�OSy��x�_�d_�F5���ɥӵ�$�6z-����)�8�M����Y�_�UH���1A>���7]p׈��m�W4���%��]������a1���S����؝n����ȭ�3@G�� ���E��r�����L��?&H�������l��c�?s ̏c�U�M�eAT��9)���]pv�N�&h�A���{`Y�G/�R������O�i�A��i�q�Sn7?��I��2s��)���HM������km�s^Y�2�˛	S-%�j�P*��Q'l�ง��!5�>uM$e3_l���&6�]���Y�^�	I�iDB@1����@�%q�N^���M)�Z-$�
��a��*�����%��w_U���'��Q趺��StZ�_����f�D��S��'���t8I�l�&ަ7C��]u�[�±�WK�ma\��bL���2#��9���rd��zU��t����G���^04Y�ܖw�io�+>:��1�h~� �d�֌'4I�����tm��+��'���9��;��k;�«�K4�/L����b�@�n�J���kC���m�<ަ �&EV#��7��{B�A�ũ-Զ�@��6��P
ZJ�/L�p��i����N��Y��1枬6hZ��1��CZ�f��i��|��b@y�"�%��j[��3_㎪��5�wǹ,FdC#g]|-d����}���S��Uc丑�Ѫ�&HE�����8&Xt+*�Tm�-�d(áE������V8\��~���yL6��W
�������W{�ߤ�q�/�T�����=��̯,�Q�m�i`4<�����{_�L� U��hqA���Y)�a뉉W�ؑ�j ]�W�y|63�� "u�,��M�0 ��G�$�^>��Z�zs�Q�s\��u�N�*X'
(Á���PD{-W�̈́�&�I��;ƭ(T �ɠ�j����JN��s�X��� |17K�B[iĥ�,�W�z�-G�׵�:�Q�K�>��	�Kޞ�t_�TWe�iKom�U�Z��Rz貏'T}<�)����{B>���ۖ���k#�"	�SY�4$t	�G�8�����G�,G&��
�ƻ����5�lMH� HEZ�����:��œ;��ѱE�1=Q�Y�Ӛ�~TPPڜ��Vh2�L���FY�"x�`R��C1E>�`�f�mO%��+9�P����uA������?��Mt[2�b�4�e�G�k�ih=�������V/�D�#`��ND�a9�� ٴ%*J����ߌ�5<����6�P<�:�R�â�;'\����`d�x��o�7&�q%����Uc<��3%*�߸
p�_�ዎ��dE�%H�=�Lx���E��i">�U	�8҄hp6�C���S�[E�v٭��>��Y�x��ۅfB�+o�l��V�
C��	#~� T��� -ѓ�Y5��|G�a6�:��7�� ߫�b�yn|�~/�j�x�����v;�����>�իO�$��&|��X%�~��aM��
�0d9Y����O�C�>
�tI�|���e��y
���wQ��J��*'�;܉b�}3鸔pҭ�=Ny1���jj��r2����f�O���Z�]�:�x�=��n�k�qw샴�k(rz�{�e��z�ήr>���=���!�o�����>��]O,z0~��r�����:Hh��ƚ,��	��o���,g៤=BI��!��Lz8�7u��&'�*�g5#x�j{��o�%v�
�\��G�*�#z�����K@6�V�
���O�¥�ˤ�j����"˞�Om`�[u~ �9)�7�y�x� S>�A�R����(�K���m}��I��AM�� 7i�yĕ��uN]� e5Թ3���j�aD>�-��֡E�e�$��
�8�c2R�Q�\>��o�~����`��#x�\�#X�l�z��(�W�f}�K�j��U�}#ܞ���BӃ��n5`��P�$ǥw����N�?�Y�����P�����l?%�e+��� co����rG7o���7��>�;5�g���[L�@L�������Y.|�S��ʯX�b��Z�F����1��-��#F�R��!�B��'�՝�gC0d�q�s�B_{��]�K	n)�6��E���R�^jQT�����KC�)�+و_֜�8'7_��� S�l��}@6|��8XiI#�s��'��y��8��m�,����&-��0�"t��%�K�:��W�DM�����r��	��]&��L�{<-/`��=�u�y�P�ͫN���B�#�o+�^_w��ϱ��RX@S �����÷��ZG���\h��~
9��{|�VDG��H��:�&\EU�:v��1J��㮻�Z�$��H�I�FB�����Vh^?���9�~��� �����B����oك�pS��G����KS�
7h�	v7�4���P7�����U4J��H�E�<���C(�)����8�SIj�o�1�u��4Mk���"�&���в��$6����p����9�}xR�a�w�dgT7�W�s�bO��<��Ư8�&�腦ai��
��p]�h��y��d@+��x����� ���.�*D'4?��Q��)E�R�F��ܺ���PMn�qPI�
ˢn���
0�'@����r;W��[�$�T�m�(�F���%~P	�/��4�9o���=�ր ҭ
XP�ٲK��ÑрN3�-iU2��e�a#h��((��7�w�:�g����%y-2^Xfu���#eIօ0�jq�Eu���cB��h�wWc� c��E���.��	w�u@�A���;�13G±���O΋"�� ���RU�й$G�2���#�7�b�{}��_%Rg����(T��~����4�S�������Q�v
�9>������w�y,ҟ� �Q��zݩ͇�Ij��L�D6�q�\0�]7��@�Zp#�sOSa��!�x��:2�ZL��az���7�|����K'!n$�&�bf���_����ε*�}I�����o�TFɗ�C�/M�I�aY\��P�S �E��^��!�/���O�%��|Œ��"t��z2ZD�,D�he6�{*�t'�Q��6.h>��`��R�z�+��{����w�(��a2�!���>D�h]�j�t�b��f�7*�&�[����j�4���E��[��MĿ����z28����Ͼg�6dl�.9����/�P*vDO�*"2�� �!B0S �Zv6���E�6��?�l�F�����j���D��KC�g:D�8�hC|}F�`(�\ُ��79$��a%�΂8�a�	�G&G$�y����+V7]N��g�e7�(��HY�~BpG�pCOBi3}A�9�jE���P��VlXW+� �|�����YF\7��2{_ϟ9(+�r�����Ayܪ�
걹����>���eB�ܲ�vK%�a�n�|���J��W,;��ΪQ���q�j�MB�ۣ��	p��n����ل5�d�n�i`�%�#X�i�je�1)�.����@��Uζ��N]0uܿ\OZ31D�f.sA�v��x�QQ&s��Y2ؚsb{��i�6�߈M�۠�%,׽l��ӣEH.��!�8)�e����`vC,���Y~��2�����39� ɀi7�0i¤a[�ڈ�����U�H&O�w��F+P�T�Jm�Rr��_�Y���ٮ>v�Z5$1Bҗ�C��}y#��g=�ɸ)�KE2J�ܩh�6\_���
�aɒ���}���8a��ꕒ?MLhl���T�'����[�7�w��	�v����Y�*�*�݈����ΖYm�O	�������Ȕy]�V�C+Ŀ���2KZ�4�nsHi����K=�X%�D���}c�=1:�����5��m{�	.�è����;�������(�,J�5�a]�#-PuX�����6XN� D��1j\Ƭ��b��I����&�-���lf��g	�E�ǀ�z����Ɓ�1Ǌ4_V[^$S�����}B"�$���7�4� ��g+�M��{�C?Qn<��2���y(��d&���k����G2�1��eEI����!�3��h4sI��dg��|[S���! ű�
�ʥ5�yG�bD��	���[�,����%o#�m��
����ga�ٓ �X��{ b�;1�Q���*���W5��jtܵ5f�}��u%��
9Z�F�ƹ�	�e��߃��Y��H��jZ�����u���[f�&v㾃�T Yѩ�=��m����t���eN\�@Q�je��5>�����f��x���Z%C�ů�����;Q5�I�o�ɒ+��.3<�x_������㹦KS��_�wW�� B��	iB7Vl������b ���z���?��e�ʯ��Fɫ(2~����3j9�����֜QQ��zrL`��\~���b=�� ���K�$=�.~�,��j���}+�Z�m	����L��1�h������Z��4fT��i2���q���qp����.�8�3&�u�"������gc�K�|Q��3���#�����"�d��g�0˘������3&�JW����èr�wj_ؑ�e'���J{���i�&D��k�Sz�O�_�diTV^>*����s�g�'E=Bi�?^d�wQ6>��gA��$hy\�B8ġY�gS5���N??��dβ�VP��s>��j\	�	� ,�vn�������_�?gsQj�s^ֈ���i�A����)��L5[�X�`�]\��p��8�e8��H��Z*c�	W�Q�#)�[���_��wӫ_΅@g@0�ٚKtr&^��*�ᗵ��M\�&&"ޅ��g��Z��>5�S����x3Q�L���Ӄ�8���5�7ږ8�h����1����+~5؎4����/0��Wz�U�H0�I�B�U�& ��6��o�H�n�x�鿪,�N�^(oZ��jyZ�d��y��I����4z�MЅwA|��hr�]���W�r���K�`�G[)>%���9TL��
��P��+�ݫ�
$�!ү��.g�I���Z��Q� �b������ß�#W2���OȜ�%T:�>�����m�U���4/A����?�y�|�yґ�X"�ֶ��N7H�)�j��1�D\��Q�!��(s�Q�&~g+g�׺�a�r�Y�*c���_�Kr�1�urS/��״dJ�Y7P{x���F���lq�yT~�a���\#��C)|m��l ���H�މ<��-@���Ӟ����H0_��㓮R�X*���'?D�]��V���υ�o�L:�e�v�����9%)���f2���vF�2r�%�廯�l�c�+�=5rԛ�M:�#�e�����ӵ��l�x��?sH���i+9$p�r�y؝���� �Y�01X���xPGm`��/x�^o(��_y�$q�Ǿ (*U���?c�T�\�#�3��a^B�:��X��՛�uCs���]�����4� ��>�;G�1�5�#!5q3�kA[̼Œ�bV���E�,ݴHT"-������g/�_���v5s��
�Ʋ�����#e̸�a��йg!�>��o�Ҕ�m���=���`�A�4�I����٥��_���X幺��-d�h�X�W�,��G�pJSŖC5�	��^I�J-�O�qz�	����\���&�ҳ��uܷ�2�@�0�7��l���ށgf(ފF�@w�Ȫ�O��O��N�����	7��^߀��J�h7sH� qHDTw��ȇh���b��d��,Ŏo;g�Bit�O֋�K_T�,�� �BlR_p]���?Ґ��Y�0S���ݼ�s�"�4��87�I�i8�s��'�7 O��G��?�ZI��*S�GNs�c�m�q�-�v*oa�7��u��G�uMU��Yr��GӤ5�X_l�)�|9�ZBMs0a*!��� ��q��R����e s�r�	l���>ed��{_?��@L��[nkz��2}�ei0�Ҝ=��O���+w�Ԫ��5�z���ǐ�;�����( W�m�r7��7R6�1��z�p��X�<.��Z��c�o�^\�xZ�E�=W&�|��T��Qީ�6�@�+Qh��n��:�+r�"s�4�8W�V�}�����M��ˈA����{���<V�4
U��&�?����˵0E�$��
x'D�m����J��'*����vq���o����:�ڱV�n>�#n�Zx��U��Va�������dv>����ٵ[k>�w�!�z��"{�E
�2������g�C!qn���K�%(��ϒ�:F��'	�F�y5�M�W��j5�`�4�f�����Y�m����Ħ��i�+7� �~�ߝR��H��d�^�[��5 �+��D���|��oO8�}H�
����*�f��"X�5V��#�9Na�~|����[�k��Y�R|k'�RWM���A��KG� ���
.
t])�����X������lf�η��&
��.)�E&�|�H1W��'h�dW��ôcn&�}1&x��&p���}�(?+�H�Y�+kq8�%�s^,�&o��L��X_�۟9�Uie� g��έ����R��%p�O}I]��#������]�:C_� ���9ur��+� J+�Z ��<��Ӓ�����}���ꆓX�O�fJ�x�n������.��K�B��h�Z�LGNO؏9����ׇ��M;�{�Y|ڌ��8���~�'R�#�3z=�F<J� x��3�ߐߑ���V�Sǧk�,�- ����Дd�%>!���s��DLQ]�--��۝�8�2���� XG���pa,�ud	W���<C���./W���_|S�i�6��?�F2�̤l>$�=N�g�:��$�BK�X��_n%�E؜"L�N����/�]~!ZV.��Yc�����BԪ��\�Vc8�]�x����'���j�m?��b�K���J�ɴ��k����]����s�_���9��W���<��Zkfq�Y�M��?�뙁�����������g��5�ۖ�n�[=�`Q�5�ڐ���␎:,���v�.qk�H:vU�m���C���s�����X#]��*r��R:}�6�F$���+R P�0p_^#Z(Ҹ�v1H��������ݏ^Uj�^2zs�a���t��d��tx��z�q!]Ӎ�O��hRI}��8Q�,W@��|#���g(;�(A9�G�+.W����뻣�0G�+g!�QB'����u	�xr*̭��.C�:C��q!gX/�0���1>�
�L�w��"��n��t@T	�F������`m6���W����;
AR�^���<c�վ�c�|�[ Q'�)�G��[_[�Qׁ����X��k]�GY��OO�E�apY�O�t�I���g��V�o������R�7-N^-��W���<����)�q=]��`�ƿ���y�sM�z-�SV�P�} $Q����A�x�G����Z�!�U5�TӲ��s1�8�ݯ��ģ�!�HꖚD�2ÀZE ����	@���;\"�U�6��D�0�ZKŻ���n�IY�/l���0�bq<l��a%�2�^:H����7�W9�<�'��E��}�Ֆ>GAF$�b1��[OM��,����d�bDN2�������!��%����ά�Lq!���@���0�Rp�dve��߳-�{J㥎��~��	3}�<�3�]���L�ky�M�:~�%:!�/�
s��ͶHn�Q��WǲEMa����P�Go�7ɶ�M$�ݩ1��t�_D01��uY��_�7��z�@���*�{��G9�@Au�J���`�S?�}��ܰ8Z��{�((�>��Ǌ�G�v{dz���>�ŬQ�Á�����`ub��bi�S|mղb>e��� K�<ȥL>�C�R*:�v[yU�y�ͨ[Z��8U�I�%�� Χ�R|�L<٫�D�+�?�d N���1e�ڊ֦��Jl#�	L��B�����X������r��@	nNP��ofs͗��}�;ڐC��Z�>h�h��M&���	[�K�8ooQ�����P���!���p�r�����׋����B�i�	=�:�.��y��ruDaHӾV�q̻�}�E�N����}{ǅ��a�'�(Y�;���q����P���+��/����Z?h�XQSPSY �B|��h>o�S ����'S�A@T (aP�l(	����e��p��٠��Պ�n�VM�,�SE�n$�}�w��{�p�p�X�����$̒�sW%Ŧq��N
ʡ{]<:y��$x��[m��U2��VĲ��<iA��\�=�!��?G!�j�T(es�f�VH��"�� �M;D�_����es�c>;c�Ki-�t�Vv�_�������:��:F�����l��3"��� Y�����j6�ݐ�x�lm���U
�׏�rFԨ��g��XҸ�kV�O�X��/��xOl �*�,302�e	9�j�Al}��R�@Q0�:ת]|�?O�tEn[��b�!���3;�/x˴ʌ���� �`�v�X�hh�'c�.$$�#_��'>!ͳ�������>u��ɢ�~�!5j]N�}�X��a\<�H�1�G�,��iZك�D���F�����Vޢ�%m�Z��&5��]��c���
7�[���?A+��,�*�w���ԝ�"�,? M���lh���/���Lś/9M�a(���w1R�����|�ٝb3��4!\qC�ݘ�����g�|�[�3&JW̚qt��ޖ$ߎ���;kD.�7��=�Yf��oM���۰�O�M~���Y;��_�?ۂ��������v�A�������q��9�E����P�U
�bP��+A�=�I:�UM�O��w�1��~S�uk�����e�	Ϩ�|�*�/BGN���� �y��pa5�����^D�O2�v�PR�2�(��:�5@b�r��A~δ�#���)�n郂��JG��pr��.��`T�5�c�2�5�i�8��S)W����F/pB��Ư��om˅Q���Hu�����{^83.��~m�� �y�ݭ�/c%=����v�t�l��_��)L��Q���ه�ҌJ�y��:6�v�]Z������(3w��h����+���y�/i�k~�bi=��v�n�q80oT��l�����Ok��W��\T�2Z�!R�Hn�2�<�����dG��,�J$@��zDX�"##Y��cé���ᑓu��d��d�5Q�
�`��y�\�(�}7��=�����ã�$%���ؔ���^���m���.�s�Y (�pR�����x�����Gb� ��IJp"�_.��VG-r��!
��B&���d�n�R� f��1,Bj�_�Pk�3Ƕ"1׿��������W�ߎ���v˫Z�/��t�!�?�Q����0���'�QưEV����k�K ���姚?��\��R�y$���WEj!����CZ�C`cg��֤Bd[?:��䒐��?�^Q����oL�0�E�p!oy���*�h@�'�ݩ dN�*ӑ*?n��o��a��v�2n����f�py�5��LZSᴘ5�g#!H{�7��������o�<%�+�}L�Ic�[/ऺc<p��씆dGMWi�-;��E^��|w!�>�?���� ���Ha|0�����b��)�4q�-��\�g]/3���A&�֖�!Įv3)Y�`��Y��|EGs0x[��ԒŖeK�:b�h��I!��>e����X�zN*�oeL�Ls8��V�.z���q�Ef ̋��Y�᪊��D�,������r������
n5�:$+�= K�f�>�[_�f���WV����z拿)Y����T
�!���]��gYt[>�I����KK���� �����j���8:��������Gg�U��O}�s?�\ٷ��ؔ7���zp5/�y�F�݃h=�@�f�
SSf�.zfޫ	7�-?�ݸt{�ʹ@8��2�e��5&�CO����
�:�^�
�+o�K�C��vq��$gk�(*t4h4����1���]@u���F�$���JW$��B۳��;�@˭V�"�46�ώPb�;���5��s���q��� )rO��Xt/�Y(a̶�˴,Ȏ?�nA���1m�Z��^'�BVO���5��=JK�u�]���g C�3r�R7��yK%Q5�0���n�_ 	��9�߫��`��~��MPv��Żڳۇj�굌5��d��P��� �[�[��u�'��"�7I{u��p�0sfaː���_�/q�!�%��,ۃ2d�>?����#X��t�g�s��N57O4Wa�oh����D����&\�\��7��	��=I�+���-;Ew���qH����-���(o�D&,-Ƿ����:D���8�C�"� ��~�����?'\*�Wņ�� �T��_X�����ژ�6s[�*&+v)�(N��A�ǒ�`�K���@��꧔��_Bh".-qD�=�K�.i,,�p���KZ��?��W�e��gT��?�6���njb4���ƙY�, D�y =Ş�(�[�|2�Hj�j.�~;����V/lc��u�Gz���^��i�T���ꮇR�w	9���4��^;����F4c�i��:���d��<O��CT�	{`
��HRϢ}��G���\�%f��0Rr֕��$������J�o&�څS�9'LT͓\��1���.�G�B�������2�d%#�~��JE']�5�I��ѻf+��HP��{����,�J�c �-g�a	&�㙇.�-A�������H�Ƣ(�����L�WnAbg�,߭�����/�:�E��a�I�ݠ,���T���./�r��_�*�Z��תȥ�%O��ӈ�*;����j}S	WXZ���Uk�S�'�g�+��;�Cr�oW
t�#/U�	�8 �@o�W[�KbP��pyPq�����xQ�d+��%f��Kl��8;��𠈫�p�sl��J_a�0nؿ2�CWg�P�kI	��?;.���6_~�ΐD������#��i�%v�A^��Xo��l�?4��3]/��x�(�Qj�F�ľ��&Ω3x�c-�y��z�$�0����W�Wg�I�>J���� ��z�oR+$���E���64����}{�8?7�?Ƙk��oG���'�TcB%�2�qG�t���d_~ǰ���&��"��F�w)_.�5��
�ٴ�a&Oma��{y����7 ��:s*ۗ� X�{U�#1)��'Hp'�����i�Q�q���W���.t�H�l٤b�(�����]�E�+�*`
�!�4�y���
�Z�I�$VÉ3\�������|�*VA�KQ̔�zt[�b%5�Z�~j�<Kq�*����!Q�W��9Z�E$��q����w�>#�|E+x�N���4;2�K���=��@�o�<~�>Ϸ����7!�X�*�{�����������M��XIE�ڬ�~��!�>�e?j"T]��h�ww���6И0��	��I&r��]��Lf�(ۑ~��[$N2��E0��.��:��gsxs�u7 �&����d��*�Et$p���?~>�3�f^` ��֛��;�6h۬NT�Z��]�:�Ր��/��e�R'd�!�)�G>�ќ�p�x	��?i��0OK��-�&���oT�=��&�1����iu�XB� ���\�ݑ����k� �T���c)�]�C^�\�R8�����RfS9�
՝�{�҄r�EWM��k-��	���+��+�l6��̥��=x�\'e�,/-�N�*(��&�v�6<��B�1]��~_��9�3�ĺ� i �n�)��OT�1�=H<C�/5��.岦����Y!2�n1�Jq9X��rڥkܩZQ:S/�Y�fc?��v�b��p�)54�O�ք_����^g��b�.͆S�%�ߕݻ+7��%cd��<߷���
���ߟP��[ੰD�~]�g�'�?�{�t�����z��nCށ֊�ywB�[v�ݨ���-=���[�5�ܛV��a���ӧv;���%�Vo�LI��iw����[5ޏ!���~��T,����f>�ږ��0��LU�8��X�f�����RZ�bm��bH-�1h���'G�����S~r�UW1mζ����� �l
1 y�hۋKH$�.�+���\��̣��Ȫ����01j4���J�dI�?���a�M"�38���k��&�u��J4~T���U��U�;�`U]�y�*u��R��h��T7��F �e�Es|�z��k��(ɝ� ���gǑ�wz����S�<�7>�v7������6	+�_M���&K�k����CP*�Iy[�-�:�*u�{���_�Ч�8}�s�U�0�W��$J�v:f������9���NM HvL��«���8�% ��vv�Ӏ<z߂Kr�y���è�9,��$����b�짃��r|HT��J��"x��i�d���S�i�<�� `Aa 3��˾���K>L�N����UW�	9Ԯ�ޞ^����=�0����5"x�gl����U�C���s��kh�ۑͯ�|��2x�!o�D�	pf�)�ߛ�<�z�T+�C��ִ����=���u���?~�	\�gA�4�m%�J��M1�
�ky�
J��)n*����1��.R��c*���U�!'~(�w��ޕYX��z���x��«��tQ����U�q+:4�/ S���m�>Jū2�l��bhI��'�Pf�g��gVg񢪵�L��6<�-��{[b}��:2�)�4��~�7ʘS��ss�t�e�ڃS*���R)>H����X�CoȒ�$vE:k�x7�d����&V�w� 0K8@c�m�wN�;����� �2�p&xqsA �d-����h��.��6��~4�b��C��}U�)����\1�vh�ҒV$Q�k����\!>F�>W�������C7eUB!״N�ڒ��h�M8PIoH2��6�GȮ�Q���G����i��ܲ狂��#���@ R�T눪^n$oR�Y�D������n������N�t��p,&Xdy%�̩��A&4%���������؍�z�訅�q$���w��N�]2xA\\�M�\u������<�@:$I�V� \���u��q/�+��:�8�4�x˓�v	�&ςz�����+�.��\[���#��Y���Ut�2��K��vX�/�xW�S%Ƨ�����x�&�ΖQy�Q-�㐷�:�\C�k��!KI���J�f2���	�c�%�YaB2m�/�z��i�|_���K�� V�t�3����B�	Z��Bi��@X�U��Ayp"�%E�TWjӠ�#R�
Z�pR����3z}��š{����a	�`���A���tS��Z�ٕ��8�jR���<���D���U%�8��&%�<���"�H��;/K�ϙ�n5�@B������%�v�3�>��\��=El�w���i�l�5�	e���8v���~�8_9	J�������+�,�BC�	)ܝ��P�(���Ĭ@��Mg-�A�=Q]�S�9NL�3v����A��ƈ9�L�y�_��4��Cm�Y�IQY�[���\�3��>��uv���o�:=txP�g�}����|���FkOn+����0٤$��*�6��Q i�R�Խ�0��(�杚-��j� E��@E��SNe�	�3Ó�
�#t��{p	����{~��C��X�K�sc�z���k>�\��W��@R-꜕@H�Mx�l��h0q5+����9��E�//J�Z���]o�d��
��1Ѩ���<'��%R�kVoڃ`෮������SE��KQ^n_-�1��Q������*DV��h��V��4���	�u�7��(6��,��Ah.e~�bm�L&���x�����Ay�&��=�㘑�#�R����֛T$R���ָ��a�&����I���� ��D�|m��00��������� {��\�Xy���0�3�$�_W���*h���.`�ndk7��B-~��7˓�*��s<��`t�7�сK��[~tG႓k澤�>�� ֚��q�t��iܗ��>�gɑx9v�I���x�0U���o�h� �Mw%v�m|	Ċw�4�w�j�;6\E���0��Q� &l�j�$�)�]�C�>�p����!�XR��Ki�m^�^�K^M��PG�r�:�f}���_�Z�O�g�0fs�ɻ��"���bH�/)O�:&a�C�Β>q�堘�k�h1wӭGX�;��X�Bě��
a�*�O�C����p49$�6#	A����=�����E$��_.=?�3W��T"{HeZ��ʠ宙 ;d�6���x��=�����K�R��#a���I�*��Cvh����CE�!�_�������}�(����9z1zZ��/�<�u4�4�yl�a����݋fu�rb�?�ׁ�����������ۏ(Aގ�W&
ځ��N����T����A���:�^s$-����G�:�%���
�/.��1>$�蝶J�jA��k|����f�	7��+�
9|�sP,��Kuͱ`p.O����j�^C�����:d$�	�H7�ќAK�\�k�V��q=��~�z�U-W�UNv�}��Qu�N�׿��s��q+bJ� ��_5^)������\�A���M/����	\o��l��RvA�b��|���٭���c9�s����R�e7LLl'��,0k��+h@�|�xb���;�<�ʍ�<��X�[�Y�v*�+��ĸwp3~���&�Ĩ>#�eՓ�<�0�Jg��Qo��Q}������4`t�y�ڦ��貗��Z��Y꥖�0G
g\7#K,�����%��~!J���+V�Z���z�2� ���0�pXo'H�?����F����u�?��8�85,�B���pv)��8��!5+�
kL_#eR`Z{+NM>Ḥ2�(<�Y��G�I�C�>*�U���b��H$��Dp�R��}4�⿂��^)'sd�E�wv����ot	"�}A�Ko<*��%v���<@m��3�Cv�m�c�:�J�GvVf��؉���;{�(���L�<mv� ��ߟ�W�D�e���掣E(Ti�%;�ʥ�:O���O'�4������wЬ�9���M�Ϯ��]W��J#����V2�92����<n�lJV�co��z(��vbg�7S<[zvbZJ���s�0�ڱ�H�Bc����6����b����n ���g�����1�n���U���R��Œg����;�LI$�k/����Y�!�CkU�%���g�`3ߡ1�@51l5�m�\W-9*^����<���CW�Xr%�>�n�KK$�.��
�!O��&7#x��=�����F_�������.�<{�������� ����8�S��.	��v��;�F�I
ۤ�BF��v���Z��CT��,��K��`S� ���ŞD��1�i�Ds��E��W5�ͥL��Q+t�� ��y�(��P���ԘF��[>��T�#��`�C�گ�M�a�|{�" Hs�����C�W~O�R�1-���5A���L��r��͎E%�:�lڼ�����<^�㽌MI�x(8x*Y+�v0ӹ��NY�直C���$[-���(C�X�����ٔ[���=�*��yR�-C���@����Q��~�y���3[�M�rQ�>A"`�V�)�]���?��dl7�q?�Y�[O�B�0�Ѯ�|���8�x�����x�=�Ɏ�������W1���y3��Qj@|��e�����®u蛷�X�Xߙ����� z$�4Oj1�� �(���S�Ɇ�� �r��k��:A6���_Nd`� ��u4��N�Q�\����|�*�-����O0,��xaL����cih�0����G4��e�u_�`�
�)D~� >��G<��Ó��F#�[���ac�2m��qp@L[�Nk�^��� ��E"�v4��ػ���2�e�m ��I;����������} ��2����G0>�lP��w�^����`ۓ���_߼��9��j,������
}_C(䄌/E��D+F�:���O�)���k����M!G�a��,[�O�6t�Nii%�>K�ĝ�?�&|��|QA�;��UV�l\S���}�M��6�d�FK�ɲhTR���
|*J9S�K��m<k}��鎥�!K�LƉ>f��G��sa�1v(�T�rɑ8j19�G9�<ox7�;�-"'��#T�Q�����:��x���iج}Q+��m��p:��ݧ�«Ϯ\21�W䢿d��`MФB�F:Ea�jSI��ͻٕϮ;뛧�dmh��N'�|t���#1!�aS
A1�4�F�b6
nV�h&�)t�
�̧��a9�c{�MӜ鏊�g5u�����W{��	`�y�=�G�*q?Fl,��+�x������cr��G��	�+�z�5K.��)_�v`��<�$r���s�c��e;�I���KGUST�ݩ$M(1�G�Ă��Z��x��5��b�����=�-��d���v�m�*O�Y_wһ L�&p��V��3��</�c��8�P����v���V�X�W��K�)>
<�=T}\���H�T �)�t�V��������!d�ݸ��S�ܗ���W���s[X����{{/Owm��q"oi\�M��>��KMXu�: 2R��{f�J*��Xwi�X9�Qix9��2T��^�(<��:ݯc�T��|�$��]߰Uූ���� n�V
�I:��;ޢM�eaO�Av�u]�Q� �&-�%�6��7�o�[�q��A��_�8LI��_�iaK�"����9k�A�m�����N���0;�"�Y��#�7��2󯋞A��\�6ex���?��O5D�[�D����%��r.��P�\�[d�&녨�yU�����T<��`\�AfFx�Iܓ"F$u؞��a����,��y��:�\$�!�;��x�F��ǺPt=����+zo��_J"�t���,_�2N�[$�G��[�:�u�m����<&�4%����kh�#j��-�J4���BFs�Yòq'�� Ӧ�p<�"|�+�2lIs{�J9�I;J�j�6�0�l� �9_ߩ��U�]O�~�>1峧,��B7�89Na�X��h[��(;�aP�IJ'R���6h2��]O�?$�)���?$}�]�CT�Q��E;c׶�9�$BK�֥�����)%g0Q�R_~mn@�Ӷ't�H"�j�끶�(�y�~B���U|�g��=�|�&�)h�t�'�]��â�|��"��ꍡe����[sv��U5�t���!��b��4��>QN|,��Po�@Qu�#+I�{f�o=��2�S@ȜF����`v�#��2$b�����cH�^���B�J�V�{���j�o\�*��q��w��Y��E"f�$Hںy�`h�t�C4�?�e%�2W�a���
���뵰꩑��4g��y��m��M�"�1�~�5G�}���>'*�* \kw��u��ؖ Z�	�4���I�����XRg�:M��?�T��Ps#(Od^-CR�����ԗʫ����L�
�|�|��>�,�֙_���(��Qw�CK� wגĆP�1�Z��񰚖������UG��OK�Q��� ��]��P#Y~��E]��b���bh[�RГ�����5h��j1]��'�D}��}��W{��tZ�O#��4Y4x`����}��r�MQ��VA�֘gL�#3���|�LS�N�L����e&�}@ڲ��6�θ���5Q�G�Q�0u��I�)q4;3"���u1���|���6X�VS��CH`澣�E R)u�߯�xԍ6��z�5���z��[�,(�'���/f��f�ٴ�[��Nr���v6|�M(,͖Fo���G=Lpv�T���m@=L���vגԏ6iK��e\a�TU:�bS���\������T��y��L)����08OKRYX0}����z	���T�a$������_$/�H��j�p�^cKu�?��Vo`@Z5�e4��ji1������Et�����I�L��C���ZS�%.��|�1�L�������2<��ߺ���Y_�ЎQί��t�_�\�w�
0~+�+��ꌣ��l9�m��$h>�5�M�P���k	ZqI�ON��J*T֡,d�Wm�b:��Rs�M@�d���	)?߄���}w	�Q-r��B�z���}�YI�w�Ub��ט��fr�c]��� �9>׻%��\"i]�DB��Y�o2�P�>#����k��;���\j>c�SW�k	���R׷I�A^���f����������ɃBg[P\���%F�I��0���1�.�Vu%sO�����]I�����Z�i�&�C�\�B��A���~��5n�gcز�\d��"��m{fxU,�&�Hwq1��%��-A}������P>s��Y�+	�i!
���!�'RI�\�q���nC��.h��ˎ$&{0�H��J����+krb��,�z& g���2���t9�Zf�RKϵ:��'V4��3�qgf��y��tt��tZacAK�]r+qf�>���f9�䖦��O�(z
�ډ|�C���b��GI�čkV�����u�i��1,V���UbZ �8���E	���>�~i�-��d��[oL#�7��&�����:��b{��}�0h���Oy||��=�_�ė���~�ĔQ�i��S0�~�N �Z9f�Ts�a���8n�� ���K�<�^Fe
�P�����iǷ���y4���L��F�����5�bb0/=y*%K7ù��t���Q��8}�dCE-eZ[��S�T��W�B犷��}tѧ�%
+�.n~!3f`�JKI�6u \J�L�pqnOQ�4�l{�b�l��>Q��+����,��|���б���`�)��a7�Vq�5��L��/��3�X��o�M3��E�.���_eT�)��O���6��/6�!����o/�j��_�&�:��|@���e&P��RI�j���<����j��^��{�z�㸷���@e8ĳL�BF��0넄�@|��SQ��׹�m�e��u@.n�ms֐�p� ��U�C��{���mB�5�+��ơ$�J�3l䜮a���y����ھ�X���h463��g�G�8FY�WlX&m1�FJ&�ŵ��UJ��&�����o{5ə�8{
N�M��>(2x)���/�7R����~�Z���������-����}ԝ���OJ��'f��o՛���%������wNch�O��y�Z���}�9_Z�4��X�^�E�G�䗖�L�J�9�v)�⁏|F�����N�s��?�����6�"��oM���פ<G���e��_��/|������rģ�l5^�������=#֋m/*`�Cp�e�Ɲ��(�:��.�^��H�[0�N�;�MojY�ڭ�<��w#G~���0�Tt�����u^U�%e7�q�f�dܱ<��[R�ˊ�[ƚ�iB�M��(�.�|�;STG�&�Y41ve�i���6.b��~\���6���ꇨZ��#�����g
�rm�ӕ8���Ӥj ���$]�a��jt�X���ς��h
�s<Ҹl��g�?Ca��m��ӄC�ѭ_��U�坜��#�:IO�X�^������/�I{E�u^æ�5A
i���WI+��n�f�s�SЁF+���q�؇نK�߫?�!�D�2�����r��t���� ~��oP��q���ՙ�g u5WbA(��b�b����g��@�柗����\?5ȑ��y����4���Du����R��3����T��f�L��z�~(�.���4-H�\-���z	�ix�I��(v:���W��� rX��B9�&�h�z�2M⏣*�o�(��{����G®2͜�E�l�=�vC:r�Z=~�	�s(-D0S⵱\Cj�VP�@VT{ōت��xa��xeS���� �T�#��)���w"���N�b#]y�ެ�n\���[=(w3�㼾E s��Z1$ �����9&�Z��{�e	�j� �yG��1a��X>Q�����jM �Q҃���=8�j���0����p9l�>˒A���f?���[ލ�ۄ�˅LEJ�XWr[�l�2��r"#�Ԉ��-��@���?.騉sˬ��h�I��WA�vC&�BL�u��N��4w����W�{n?(x��S*��$���`P�j���-�������4�S��b��vd����3�lB]Dh��� ��P���tCP�6D����zf�;�WƓj��i�c�*ϗ��S��r����}��3W���UQ��-	��U�+k�;�̝}|���5}=6���S�M�� /2>fI���,JBi�g�T�MӀ����z����Bʷ/ؚ Fґ:�?!Ec�K��
�`�%
 ���y�y����
��`E��}h{@�R��IE�ƫw��u�q��bvG�<��N���!��?|����'�JW�Z�tV�q�$E�T��쿸�F.��ް��s��?������nN\�N�>�'!�:(E�0�~�P�5��EYn���7f�eARZI�aF�:[��� (b�%�o
^����'Do���DG��>,�S��R���\�d��A��R�o��t�!��O���\�g:i��'i��I2U�0��K�k�TO�����R1�����p^���@>�ײA�\u��ɽ�N���!7�cn'y��.s�yMK��Ӊ�n�����i뢧��(d��8��r�y�1Yփ��گ����)f�?�K	�I���j��׍הs����P����L�H^����1�ڥƔ�J9�`O��e�y��͏��ꡩ�3�I9�~+�'A������kp
�eF}쇐�`�h!Y�d���9���t�6��	qGWq�(���5&���1����*N�3w>���6���[�+����@T@�)�q�'Q�B�|�a�E\��G�T�(V	<H `���z��w,�q>d��ɺIn52��c��v<d�)ꛘ�)���Ӈ��B���șkX%<�S�}��Գ�C��A������rK�����V���B� e��7��}����Hi�+'�;ً��7������U�F=)7]�E���R5�i�6�o~���ļU��/3�+���{����j5�c���w?߆������1e�uXɩD����n�����e�k���~��[���]��W�3�\�&��]�,2|��j�>r*lt��7ɠ.
���w����/�Ї��R^�{TZ@u,��6��Ԇg��iً�I'��2����fh�H�c�7��M�/�vmXgzX���*��
�����'��U9�B�ϗ� @�b�T6��M�W�Q�/+h������P������]a���d���X�$�cZ%Qp�[
�/Gܦ��D���C@�s���������N���	�%��~|�7~���o���p~���/B�-�ȝ�ϱ-������6�L�F�;7=Ww���Y��We�j�QM��(+�!kL���#��u9;�j�s�����8s�!<��+��}#�%4\�w��������.(S:��|,��'��V����4��&юr��-�)dOu�:��D�I�ݭ�
8�7��̊���ԕ�_�;򺭇��-��(�g�tҭ���؄S�t t'
�ț�ed�?�X�߅U��%S;��Br��(������
7PO'���[/�*_0��'��s�{���>{�h����N^�m�$�mVSDU����뽞u��d�V�|��3�%���@�q�b�rmHW�tȐ h�8���ɇ��H
�&[�+ZٮXf�v�p�?��}��ѡ�Xp|s)j��C+AN���&�ɼS�L�M�h�F�>)���!Z��I��}W�`�K�fLHjR�=�(>�)��m�!;+5��'m(5��w�4Y ��1����J�ye4�v,���ՉI��rb�Y:����Aȶ�Wq6���k<* @Y���������`�����E�F��4X����ܟi$��qK��8����<w	��K�G�K���T�)�g>�m3<"��������~����lR=0"�Hǂ#�MO��|����O����o��i����?�	�g�+_�����r��������*z���F?ݑ>fW�`ݶ}�&�og���\캧T'Q��mp��R��X�1vvO����v2:7��p�I>��K;�\J���ض��%dҋ6!���J�4vE%�2����&x[��)`ϵKM����VS�R��P�n?z�RBX�A"�!�y�/���pe	Zf^|�(�)&����	��j0� [�dG���O9�%�*q{H�V��g'6X'59��r��Z2�أl�7��� ,XU��N�Դ�L��:�Ӏ�s�$R���YF�Soo�������n���mTLFe���u8>x�����_�?��l�Ev��������Q�?L��ӱo�'A�m�9�&� ��g��e��l}��˝Pߗ���e\�_>j�`��|��f�3�*��`!��I�D�GV���gf"S�d��L:�;�wS-P-��E����u�P��u�!��$��ӎ��
�S�`�ѓ�����+@/��\O�����;L�ޗKk�LA*�t�ˀ 6*{G:�� ��r�0�\5}V�s���{R�'��.�c���W�+&P����b��+-��Q�?W�ij�[@@�����S"X�މ1�&'�S��7=���s���eh��>����LZ���z��n�5��9�J�Ҵ��gI"Oס	�����-�%��g���"o�/�}Q�y��{-Sm����ye�}��^!����=��2�m�rTjX���t��G�MJl;�"����@��[=���!s�s�&YQU/���M�=[���������8���F��Ѐ��cFy�!'��Ps�����_���W��k4�m��e��wn^�8�%�H�?����F0����ѡ v���:��q�u�%��Gȵt�Ȳ��_L���Ѡ��	��m_��j3��|N�1V��F�W�%��{��u�b��L��6�ｎ_i��#���,>%ڧ,�}�W�ݷ�o��nb� [�~{��"谂_��pK���RZ�*m��K�	>�c����͠�:w�@>�3_����rZ���L�/�D\���S(�ۋ�H6[ɱL�ʾ�3v�3qni^���SB"0e��(���v��2d{aC����_�K�	]xI������5�f[{t��>Oc^�`5�ʉ���xDn�d��}�5u�7]{x,�&�ńo_@ʠ���d��D���N��z �<�Zӗ@���|����%��K�6"�a��A����ن�'G1o�:2F���[�׀A�,��a'+��P2�+��WP��k�����d���1ES�4��1=�5sX� �0��4S#s��af����4� ����@�O�`�hv�P_$&��'^n�y�A i!>M�6���4�E��z��Y�c|�w�g��J�Цh�*����"1?�iv�5����yEdl'B�q��ȉ�ѿB�yr	j'�zt����۱O��;��:�M�(EW��TZ^�{�ewW5���W,��`t��MF��=-��^�V���i	e�R%�$�t�w��������3�*e��ڪ3ѠZ��bxe�ȘH��
�l:�q�9r	�4~<l�/�b��ٔl�J�6�T�n�Vۍ����L�!Ի�:����� �@��|(��%o`�%����X�Jƶ3����Ex�k�8W���F����9�M�VԩCb�z��Λ��<(�f,$�
�/�K��;��@�#t)��#l�k�n�95#���I}�;���L0���Mu�:���)Ka���ü�$���B�ԡ~T���{=��ʓC��ZN]|�Vv��
ՠ]%�Ѻc��@�WVa�9��Gksd���n�N_Hۮ�q���T$��Z㡜2�ŉ0�6��r�����$����S:lxי�/$����p8������ց�)�"c�+	T�	z�V�0j��3:!44��EP��#�Q[����T+�B���zvBy%�O(���ES�7����}��[\�/�Q[��o���aS�I�V��P�+�,�^��j�8	�S���e'fiS
/��Q�]!'}��ڇ��P��ۢ�+>����ť�ˮ����K�U���9)L��h�';�����u59��9��k��=a��0�i��ѣ��I$3�y��tV�~��^�9S�[�!�-1n�y�kk̯ʌ
�n0C�	#�9Y&u�hɶ��#Z�H 
A����)�������s$g��
�4�߄��		�oaQBg
�[�:��f�$��Ȓ{;�����iP+Etl$
|~����]G���%�Nh��FS��� I��(K�m>�
�ٞ,LĞ�c��"���R���:Y�N�{̣e�%���%�E>?�g�۟?��
�������d#�B�}���
d�.�"c˴X_o���^ڝ^[���&H�U�,Q`�1b��S!�
�L��\y">��G?��;
ߑ�0����^����Br(�5މ���D40q�h��}zu�hi�{�6b� s�5�󓄃�Vװ� 8���>�3���>�����9�����\<��U���ϽZY�d���W&��\d����.�����*�K��%d��o/�GDmJLhY7=���Б4��E �4�1D/���\"nC���S�\���3���m�̽�H���-y�ބ��-Z�걄[�z`f)���V����Fc��#�{
��+S�Ӈ7��o�[8��m����>���2	X�d{2��P������X�g���
�txan��U/1�/�@�_�FgY�:�����jfM����>v��F(F壖ϳ��~��_T�z������4g�!*N��,�`�Ӧʧ;+����1��X��ʎ�S�z6����nJ��^2�&�p4�����)���DT�Yx��{�.�a���<
��V�����2aG�p�3�Źc�@�?�ט����vaHo�Y��STx�u�y��=כ&��%7�����Wl���f�"\gd�p��~Tʠ"DR�@��j+6�=!�BT�4Ȅm��uM�ƕ:��n�\����e#�^��/�y��߁[D�L:���,��>���͙�ݙ�����#�,%W�dd3�����W���u��/(��lGv����V����|����.���?nY��ߧ�E]��! >g ��SK,�{kJm�Wl]�%�۞�R�W�Qj�:��h�Z��c�; �z�E��v�&�1/}��� 7��m�&IP��:�<�,͈�ar�������ą�k�yE9�G���πE��5��z��}�D�l����^�����ш��?jϞPF�*�u8�+�X�(�V��p����?��HZcq� xΫ�R5@j�
�:^f�F"�uS�f��6�7�/:���\e��T���@��L�׽"��I�]w%��z�Sdn�s�I쀦��ɂ�ߣf�������%ߋȰ���&[��k�� �Z.x��^D~��Q0E�bk�) ���j��O�y�6{�'ț�Nh�Zj�i�+�7ӂ���2���zM:e��
LF�W޵e
��n��^ʙ�q+n�jl�q���S���N�v�m��}׿H>ԃ!�JV�����;�4|}�J��KM��HRXb����M�5̨؈ط�U����A�ǻq��2�j	s���)����Tƙ�"�L���\Ǵͮ�0ى����i��_���J�aWqjOq�R{�IȮ&���V����G�p��ǎ��Z\��e6O�d�k/���W�ӱ�4aE�A�J.�T����;�{�;Ӥp�5���4����i�Н�#H��g����h����K	�њU|��p��%��&\���xNqI��YTn�j4o2N^
���o�����`�$(z�>l�C�kd5�>� �og
�ο4v�B�]�3�PU�@P��p!��e;�zo�ǂj�fZ_mv�#}A_U����jI�t������!Z[MG��D����)-\M�rw��;@�-����[�\U�J�-4�W���P�	k&�mp��BvW�}A����q.�-9
6ћm¡�����喩	�wuG�m�A�oܨB!�1[����m���Ď� p16�������~������~��t��u��%Z/���:�a*AJZ��P��I~��m�l��DG!>��7�{��S��d
����*�N* <z �7�(';����
v,�b�J�H�x9��:����}xMh��%�N� sz|�u��'Ǩd���E��}?�����R+{�% ���w������z�b����	�K��StH����MŔ�YЫ���#)�h���Q&��eH3�ؓZ?��{����)�Qc�[H�����О>��۩��@�ѻ�Yv���h�?y%z9�O�D�ƒk	�.%
���d��Z���?��6��Կ��1Fv^o�㑧��sM6B�i�l�۪�}�=ger$�w���}����0:f�<�>9���`�="�G;Uc���ğU1AM|��n{�aFrF����������<*����I������@�s��i�q~���r�tHCɿ]��hɦ�ΞN�̮��B{Ȼ��Yb&�����邖�Q�,�3�p�ۦ���\��=���@rw^y�|(J�.��Z���|��/�	���	�D�יŖ�#�eo��_��)�Ct�j�%2�n�=-Dʍ�=]�k��T���Qƃ�?9�|���3�M��Y��M��(��� NJ`���L�o�^�&��r(�Q�����w�·�>5}Q��+�&8/�J��5��E��3�����5!7kD���J~nY!���Q��]-Yğ�9��IZ0^c�E�x�A�2O6��E�-E^q��c������`.t�.jT�7�z|�O�u�9N�4=�| kR�Hp5-^��lV���c�����89RU �α����F�Ȥ��$�lZJR\"�F�$���t3�&�;0�/���
�P�uc��J���H�K�I\jg#G���˲ی?���?��_��9h����ՁM�C�7eh��[��$vJ�
�����0{'��u5f-�e�c�`��J���0�L�M��`�Uc���Pab[�/}`��r���=$m1פ�����š3H��l´�rp9&{��QC�]�}�s4� k��W��j�;ڰee�9���wŊ2���s�k��.�V��{m�MRС�8]���5�ڹ�:fq�J�9��m]""r/����WZ%9UL>�&5���b��:�լ�d!W�z#6��d���T:��`#�ֳ�l�����9��gC���KE
�4�rc�a�ݛ�˛�/i 0N�*Ǥ�jc-|��V� 3n"��}�á\��*������h�Ѳ��*˼�bu �LAs<c�&b��CM�������X��o�φu������[>��І@f
�x�p�n���{L߸ꃇ{�q��y��+�p�oH�:h�+F:ڃcNN�Z�&�l&�}w�ٮB�&��h�%�VE���N��G R�|�b�b���,,Wb��̣���nv���������v`>M	���D�j�G����_bC��?��_���U���|+3+�fA(�1}dw"���������٦�J�,MPش��H$ʕ������=G�:��,	�˨���}��!~Oin�N����Hm�H�1*B��g&��q6[x�O�y:�yF�L��-�̞`Ꟙ��o��ϔU���o��>�\,\��ˊ�t� �A��<ع��&������d������v����D�ULWS��# �/ҧ��0�ԹĞ �Z5rY�>���+��N0��X풍�I����1@"�_>����d�Y����o�a��w�j�H�W�wUפ�}c�5͝2�E�Ir�wa_=��ۤkH4��C[>'Â��%��nw���6�$�ë5+ns!&;�z�Q�����������w�!�(�O��z�S!4w�v5�ޟ1��9���)��\\�d;����W}�
1�bs��3�X6��4
ĲKj�[:֭׵"0����cN���,�]f�E�ED'4�4�"�+�w�qSd9\�A��R�9dS�z�\�'O~j�i�� �Ȇ�� }�܄0��V��	z�ֲ�N7�P��s�G�c,��A_;�{]��~	��,=�B	�mA���MϬ�O}VM��V�k��4Y�=ן�V�o�i5�_KR�+/y�g�z���PzĐǣ����c��hǂq�6�Q����JQº�N���V�<�J�;�&�-w�`���L�2N�_O0����ٿ��Q�M�3!h����{��wO�d���i�?g�t��~�J�ZO�.�k?߮�x��2s(	�yqu}�*���{�j����Yq�^)�C��\��Q����P�H�~b�&���ܹ>�6�ya.�gOlj�8�U�0+����[)�/:��#��-��h����2�s:���xUˤwю%N0)���0p���'��Z��!�s"�M��2���X<3��y��]���<�`�MrH��Ct`f�6ҍlo/��|��F������p𑭈}D��! �Y2Z��0"+�s�ΙB��	�2�ݵ���H�]������ot�OF��,	��Sؙ��G.�<%��`��n]z޷u�1L6;�p׫�in��������ja��eX���u�n�. CY�X.F~0Y��#�t/���T�\���R��{�K*(��	��ʲ���u@�e����=��ی�?��������=�)��.�^
�~��̽��I��x�p�/�Z���ۂ��%]���� ?��$�ib�TG3��&�l����j�(]<gr��B��Z��[s�+�Ȯ���vO��u"H"u���0fL��a03P2z��&�#�ὧ��4Zޟ<�~ m�H9��g�\¶]�5�->\Γz;�a}'�x}�K�)��5x7m1ɨX`�)�A��AS�\l�<"]D];�~�xT��Q@��ZC�������8�jO�3�+4�'�����*뼒�����
�?�۵�@=.�t\́�	 �ԛh��w`F����S����#��ё�������f	ȅ��Z׹r_SL fhA�+nț,Qvy2P���,��_�q��r5���Dr���t;Q�� 8�"�4��es�:��y��Ljt���;��[�j��;���j�и@��@v�P�[�/�M��;3h�|�k���4#ʲ�"O�4j�=C��8�����M+.�Ld�'1:s�Bv�&A_�Ҡa���p؆�SW԰�C{���<�4�*�R��b-�QM�Pˡ�K�ٗ�?�u�a�2��#��ZV�6�/���[�F�qѹ�ɩ�@6x��41*�4�8��p�FXp"�;����9�6�Fg����@��򍉖��D#���M��BV0���A��y���b����p��(^(W�Dj��|�c�&��~sB��K*�:���QN��������d������	�%˾X�a�C��7-s��J��"z�v&�\#�%m�#��/���߅��<T؉JN�Tֶe���U��T�oe��1N�2vh�#��� ��hm^й��I�ZYu^�H�0�B��*�����t\+�6�F ,��ѽyN���ta�W{��$��1Q5��k[�(�^ ⪹���J]�`r4�	@'ʸa|Uj+V$�a2qJ��L���/��F��H�o�s��n��G]zD��Lp0����!}���"�^#�a��obs�ϛ4��h�����9κ3���<�P[��>I�?�yK��4=������&x��s���fJ���Qv����0���<RPi�������>��{/����kPSf�>m�r���-'�x
�BC�W}z�i�LT�/16W�*�?��Y,�ފ�󮢭{��&���$�B�j�p��*b߃������ �ŝ�Q|�?�	�ȅآrZ��w�jO=F�z"нXd�;ݶ�8q��<\ǂ4m['91<��+*`�X����0q��0��١}"�.;�	l�w�aӫ%���"t��=�M�E�n�ԃ.�A�Z*AB5(��@�%�L�ڥs8!v�zvÏL0ѻ
��2���V����8�'��7��#�����[֍�t��!�>�"��hiT��� u���+i8����� 1'�8�/�Hi�HJ����s��;�A1�ic����b 咊�3;���al�$�*dJ����O��r޵OY@h��7 *L��w�k����2V���/�Hs�[%^�^W%��_y$V��� dOJѧ�+�Z���a'���0
Ͻ\BM"D:�Wb�\�_ME�\�I�b������b@2�޹��
P%
9U�5OR�� V���A��3�����a��I�:6�Jr2���W��/Ry��b��Zi��8I3�X��P�蓋����Ie��I�po���d ω���6k�;O?b
*�vF�|�v��ً=z�T��xc�v�|Q���������Z�q���6�{���0�<�y�1���k����|{�+n�>�pら!×�����NԬ�+�Ǵ	/߅�O�O��A��|3c:�� �Н���m�ԞOM(,`�kK��6��)/i��àhR��-��u��v�$�;�t9Ұ�ǂjTM�%??����P���ș]�/��c��)�ߎf�$%2F�b�Y��8�xNL9����i�U���S������YM�L��m����K�<����_��CR�DK��.����$��S��c�ƣ�Sɪ��4��y�$h"R9�ב�R?�;�����[���!}�9&gN��@]�^_��7}�9��ϔj��h�V�\�O/��:�u?F:�w��4�*�2�����LRw�1�W��z��p��^uѺh8nԲi+�,&k���{�g�=5�{���h:��U���bT���q���U�['J���&�s�!��~Br�:����R� ��2A>��Ho�+�]�ż��k <k����&ڃzAr��S��PE�V���"0:�T����/W�f��6���S}���+|¢�k�<.���2*C��g���)�O�4����wG���0CM6�&B�_�H�5ќ.�r�&U�6�XLm ������5ӵT��[P�g'��Ի4���`J/�t���BKa"Nbr�A�x��|��f��z��l gY*�H�/<~>�%5��Q��uT�Un�j��pI2��2�2�#�O��&�
~E��{�������1Z%���C�]�/5[C�q9�_���}���Zt,��er�-3B�G�ʰ�O�*���vV/+6q��҅d-���<����7�,Ν!wmjk4��j�};�$�����N�+Cv)��x�o��	I�B]���FC%����B�gaȦm�8xWPk	�(���ۣ����(�����eM/sق���XLh��`,SJu~�փ���X�#�O��x�#�6��t�Ny�tfF��0��vd܎� Ѐ�6!�e1ּ�� C$�(������g̪��WF����Ŕj�O$�a�(�ɶ�dYymf5l%����-�(a�$�ׯ�c�S�s�%`�g�����q�>w��z��i��9@���y�n��%=܃����*aI<8z������N@���֍q����t�O*
�$����0ü!���@�'_YQ�v( Ia&��̕(���.�s�t�+��Z�b�{
�褕�����/h!3���@���Q�$?�N8dS��G�S��ڒ�2#Q'��IZg�F��0/�G����>�g�Qk�m��G�=��Qnӎo��G�8�I�5���D�SS~_)�E���ѣ6r5!��&�Zw�r�X�D���t�S��b�	��}A��q����ijxp������l� rY��<|�u��^�3 ���Ձ�J�=vA�(����F�U?Ie�[Sߞ��w_�"����i�Uc�.jA|m#����_���+��m�妑E+��&����q��G�|�Ț�T���!��Z��^r�*�޽y���|������:��(^T�IY��]�M�:����_��<�JSu`%��*� OS�����oŋ1R��t�[9P'Mx|��&(|uK>����z�H�o�O�'_&h�� %��M�}n��I�����hc�|u#�]��K�"(5�ZP��Hx�@�<�fۢw�;ܨ�p 4��6�qK��T��Ѿ��jK:�^l�Ы�q���g[�S�ŋ�����-�W�%�"r�kZw8-�O�⑈>��S�L��x�*����?���� 9d���j8�S��sϫ���Z�i(����uƹ?	�#R�7�"��W�*oҪ��aݏ`���$�X�X��5C��8�e1%YJ���iFyۋ���C��9�-�$'j���s�k�о�&}��;�*7
�wo�M�R����*(z؅�FW5`�O�<毶����ίs��<��ԊcY9Q�Eq'�����dX��	�9X�ؽ�v�-kL�s�Ʊ�~nh�,��� �*�І��P{��I�dG�D��X�焳* �/��$ֽ�F��nP�>���?�_V��چ�?u�}r��s�K��N1Y��vX��0�:p�%LQ&Z\�'����E�E�����a�|�����J�W���vPO��厲���`� %U��.o� ���Z��ݝ�ғ3��T��&_����.�rAQ6����\F9�$�P���:�[���۾&���� q+xyRl~�rX���R���K3<�I���p��(.�_߰5X��~lO��D���j�T%�6~!�7N����m�U-��3�h(#����{��f��R�Jj�<���g���^&��?>V�4=���a:���2���{(Q����1��u0i��; �H@��]O��$��EW,H�!o�-�ܧ�zb��t�,����}vn���-�r%�>�"�V�^�ߞ�ٽJ\D�O�^!�[~`l��V��*ޯ��mM�	~Φ�!���)�ܥ��<?�a	4��,+���8R6��q$a�עx.��=��|>V�5��F,��>{��8���Ǉ$>s^��8s��f6��z�]�8f�7�E�DU��)eי�@$�r�r�jtHk���lL��;f�O4̦�NOwUtՆ�m�Ӎ�㤍�9�Ŷ���Z&O6�����޹�*����Ng�@����E�y�]ۓ�1��x����RS`9;̣�{�9�f X
�\�~���|s(�#�UH�=_�����sySj�^e`"{��1a���b��=�-Wf0�C\.�w�5?����sI���I��J��O��wlB�-�}/�On�N��{5߰_v���nr�&��Av���hۏo�ol])�@f�7�}��
�3��T3ܛ��EM������Y%�6x/wX-�5h�NA�/�2�T�/E�ЀF�
���7�{;��� �aQ��������H-̀g�3����?�IW�'F�T��[��X�zGC]����H�ȫFƭA^�R�
�|���������/��L�Z	7ϴ֓v�'a� +��"���N�|e�Ԟ>�o<���=]��e����7��`�\-<��������5(���S[�|H2�	�A�g�TX����b�nۘg
�2�?梩� H�{USԙ���L>����kW��Nt�jC���V�-	כ)s���f�֛X�DE��'�tAb�P:��6+��W��"s����g%����j�"��BO����O,�|����k<�hL�PK���~1\��߾���D�����_��
@���<#CU
���	�\�t����K��3�Ʋ���i�j\ۋ�zT� >4���{T�f<��凎���{��`i
�I�1f�j!)���h����$��I���G?sBsE�gެ�X�,�L��2A`�����kAH<TPI��h�۩ �,n��C#��S+����a��o��^uV��m�=��=^~��l��C�8����(浓�.�P4maj�ٮ���_!B��i�$��sg���Ҷ�J��E�Bm�F|)��F�?n�Y � [��%�̛
b���I�@��>���grq̶t��<ƽ���Ɓ[L���lk�I�90���U��=��,���@c []Y��w5���>�����:��^.��_,$�4��/����,/iq5׎��Z5�6���%򌵼T&�&�퉜��,�Ҧ�&�}��l@;ˀ�j�� �������m+U�̀)�_2�����Gҫ�q[T��^�ƭ��*^Xi˳����דr�;c�.	��ַ�W7ڧ��h�k���IM`^!��&��������R�Ba�)u���s�/�����*K�Xܺ��A5�$�n	ї�lN��ZD�yYnS����=/�5z�;+���Us^��m�lk��J���H�qRq��	p_����{�O�6P�IԬ��xA<m͑���Pb��`˃���c�Q��m��+�����W_i�z�`7�t�.�oX�Y�3�j\�U��A�a�o���h��,eKAVlaK�/�ba˔v���q½��S�-<y�s}C ����2�p�Ӑ�����/N����3�C���,�0u+6�U�y�����ᾔ�E�*(���"�$K^5�
W���"IM�p���c/ kk���}����)�AAg����.0�XG��jV
4n95�<1�N�=�oe(�|s�7���G��L6���Æ_6awވ7�h����S��k��+~��Q�*�W���s,>���̥T� ��d7�L�쮇�4�bs��dN�{[�5W(�4%�s�ɒ�Z{�L�0�;<ɨ�n%��k�jֈ6�]?Ls�?ߢ|wGuê�����_y��Yܲ��婕 K���-��FA�\���PT�<K0Z w˪���.H��D�}+��V�I�f��������G���:�P����v�2��r��j�ޢ)|M�:����u����_�EV��9�E���Bgqpdb��t�5oc���vZ�� J����gKC���8��8� (B�[F��WQ�z@��%;�����+�=[���E.,�(8���0�����E�y\C��@����@�:dC�K����:��X4ٕ�g�E����la0TmF1�F�����O?QP��j�Y��QrW��I�T�P���dʧ!�����^��p�D�%�#йVFT��: �xr���]��l�x��,� ��!{*��'��a/a��m���m��78��=�Öq:�<��cAzg7�oό�Niw&kR���7
�Ň;�27��Z'�,
����h����~,7��q�A��zD�ddJ�b�-2�d��~�W�l��.V6�#( v�θG��FSwD�x���� ���n�|�$�M�x���K�N����9 �1S�(iX��]�)G�:y�^����S+dH>�ՠ���V!R���7'7����p�R"	����D����n�-��//�H��T�z������=�ˋ}�滛F���[;�p�+	8c?\N_�KƋ���m�^���5A:kR@�}��ȁCD���b�A�ٍ=̺{���\�Ǉ��_�N��� x��0k�bF̾�!����H8A����zp��t���+%^���qbo/W��� �cE9���@�C�p�3��XaYVj�<)�H0��<Uv5����mM�5)�W-Rh�9����)���� �!;s����ǖ���M�Gh��(��װih��H�)�7z�0�f��i���B]�rD����?S��:����J����;P��y=G�A���4�`�!	�h�B��3(+Ҹ^[o��E��uNW^�r�z/���ec�b:U�	G� �K�D�\H�Bv����R�)6O3���#�=uS3+��ĝ�On�zR��E��6���g�d�����G�7b�������}���l(|¡���G�ry=YU�Q�i��HCr��l�[PY�}{�!K)�)ܦG��|o��j&��{��謜���|1�3 v�=�.�IR�%2l���,�F zU�ܽu��ξ �J��[w�ƥ���x0�T�KD��y[�O���� �����+駓�WGf�|��1���V~��M�����Αm	R�;�rZ�汐��2r�� e+}��1�d��D�1��ˆ�9h��x�U�2`�̤��|c=���=tafEU�H1 �K��0X�OÒ��P�����]�T�|6��r���s{�f�.�3���HlO/��8w��}/H���S"T��jF%W����e�����&���c��w�}�ؽ��|���l̑�-�������~o{W��q�8@�?�.�G<
E���Йa!/>�cU����_���>б9�������@MoX9�Y�3HD+Tcgn�p��;���\	5\q�K3�ZjN��fxv��a