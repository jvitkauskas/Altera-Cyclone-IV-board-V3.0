/*******************************************************************
**���ǵ�FPGA������
**��վ��www.OurFPGA.com
**�Ա���OurFPGA.taobao.com
**����: OurFPGA@gmail.com
**��ӭ��ҵ�½��վ������FPGA�����Ӽ������ۣ����������Ƶ�̳̼�����
*****************�ļ���Ϣ********************************************
**�������ڣ�   2011.06.01
**�汾�ţ�     version 1.0
**����������   �����(���������Ե�λ�Ľ�λ������1λ�����������)
********************************************************************/

module half_adder(A,B,S,CO);
	input A,B;
	output S,CO;
     assign	S=A^B;  //���
	assign   CO=A&B;//ֱ�Ӹ�ֵ����
	
endmodule
	