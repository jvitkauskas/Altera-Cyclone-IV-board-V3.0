/*******************************************************************
**���ǵ�FPGA������
**��վ��www.OurFPGA.com
**�Ա���OurFPGA.taobao.com
**����: OurFPGA@gmail.com
**��ӭ��ҵ�½��վ������FPGA�����Ӽ������ۣ����������Ƶ�̳̼�����
*****************�ļ���Ϣ*********************************************
**�������ڣ�   2011.06.07
**�汾�ţ�     version 1.0
**����������   led������ʵ��  ����ȫ��4��led
**********************************************************************/

module led1(led);
	output[3:0] led;
	  assign led=8'b0000; //����ȫ��4��led
	
                          //ʹ��������ֵ���assignʵ��
endmodule


