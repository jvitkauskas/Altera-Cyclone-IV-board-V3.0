/*******************************************************************
**���ǵ�FPGA������
**��վ��www.OurFPGA.com
**�Ա���OurFPGA.taobao.com
**����: OurFPGA@gmail.com
**��ӭ���ҵ�½��վ������FPGA�����Ӽ������ۣ�����������Ƶ�̳̼�����
*****************�ļ���Ϣ********************************************
**�������ڣ�   2011.06.01
**�汾�ţ�     version 1.0
**����������   2-4������
********************************************************************/

module my_decode(I,E,Y);
input [1:0] I;
input E;
output [3:0]Y;
reg [3:0]Y;  //�Ĵ�������
always@(I,E)//�κ�һ���仯��ִ�У������߼�
	begin
		if(E)  Y=4'b1111;//��ʹ��Ϊ1��ʱ������1111
         	else
         			case(I)
         			2'b00:  Y=4'b1110;//��Ϊ0����Ϊ1110
         			2'b01:  Y=4'b1101;//��Ϊ1����Ϊ1101
         			2'b10:  Y=4'b1011;//��Ϊ2����Ϊ1011
         			2'b11:  Y=4'b0111;//��Ϊ3����Ϊ0111
         			default:Y=4'b1111;
                  endcase
      end
 endmodule         		