/*******************************************************************
**���ǵ�FPGA������
**��վ��www.OurFPGA.com
**�Ա���OurFPGA.taobao.com
**����: OurFPGA@gmail.com
**��ӭ��ҵ�½��վ������FPGA�����Ӽ������ۣ����������Ƶ�̳̼�����
*****************�ļ���Ϣ********************************************
**�������ڣ�   2011.06.01
**�汾�ţ�     version 1.0
**����������    2ѡһ����ѡ����
********************************************************************/

module my_mux(A,B,sel,L);
	input A,B,sel;
	output L;
 
 	assign L= sel?B:A;//selΪ��,��B��ֵ��Ϊ���ʽֵ,selΪ��,��A��ֵ��Ϊȫ���ʽ��ֵ

endmodule
